module Reservation_Station(
  input          clock,
  input          reset,
  input          io_i_dispatch_packs_0_valid,
  input  [31:0]  io_i_dispatch_packs_0_pc,
  input  [31:0]  io_i_dispatch_packs_0_inst,
  input  [6:0]   io_i_dispatch_packs_0_func_code,
  input          io_i_dispatch_packs_0_branch_predict_pack_valid,
  input  [63:0]  io_i_dispatch_packs_0_branch_predict_pack_target,
  input  [3:0]   io_i_dispatch_packs_0_branch_predict_pack_branch_type,
  input          io_i_dispatch_packs_0_branch_predict_pack_select,
  input          io_i_dispatch_packs_0_branch_predict_pack_taken,
  input  [6:0]   io_i_dispatch_packs_0_phy_dst,
  input  [6:0]   io_i_dispatch_packs_0_stale_dst,
  input  [4:0]   io_i_dispatch_packs_0_arch_dst,
  input  [2:0]   io_i_dispatch_packs_0_inst_type,
  input          io_i_dispatch_packs_0_regWen,
  input          io_i_dispatch_packs_0_src1_valid,
  input  [6:0]   io_i_dispatch_packs_0_phy_rs1,
  input  [4:0]   io_i_dispatch_packs_0_arch_rs1,
  input          io_i_dispatch_packs_0_src2_valid,
  input  [6:0]   io_i_dispatch_packs_0_phy_rs2,
  input  [4:0]   io_i_dispatch_packs_0_arch_rs2,
  input  [6:0]   io_i_dispatch_packs_0_rob_idx,
  input  [63:0]  io_i_dispatch_packs_0_imm,
  input  [63:0]  io_i_dispatch_packs_0_src1_value,
  input  [63:0]  io_i_dispatch_packs_0_src2_value,
  input  [2:0]   io_i_dispatch_packs_0_op1_sel,
  input  [2:0]   io_i_dispatch_packs_0_op2_sel,
  input  [4:0]   io_i_dispatch_packs_0_alu_sel,
  input  [3:0]   io_i_dispatch_packs_0_branch_type,
  input  [1:0]   io_i_dispatch_packs_0_mem_type,
  input          io_i_dispatch_packs_1_valid,
  input  [31:0]  io_i_dispatch_packs_1_pc,
  input  [31:0]  io_i_dispatch_packs_1_inst,
  input  [6:0]   io_i_dispatch_packs_1_func_code,
  input          io_i_dispatch_packs_1_branch_predict_pack_valid,
  input  [63:0]  io_i_dispatch_packs_1_branch_predict_pack_target,
  input  [3:0]   io_i_dispatch_packs_1_branch_predict_pack_branch_type,
  input          io_i_dispatch_packs_1_branch_predict_pack_select,
  input          io_i_dispatch_packs_1_branch_predict_pack_taken,
  input  [6:0]   io_i_dispatch_packs_1_phy_dst,
  input  [6:0]   io_i_dispatch_packs_1_stale_dst,
  input  [4:0]   io_i_dispatch_packs_1_arch_dst,
  input  [2:0]   io_i_dispatch_packs_1_inst_type,
  input          io_i_dispatch_packs_1_regWen,
  input          io_i_dispatch_packs_1_src1_valid,
  input  [6:0]   io_i_dispatch_packs_1_phy_rs1,
  input  [4:0]   io_i_dispatch_packs_1_arch_rs1,
  input          io_i_dispatch_packs_1_src2_valid,
  input  [6:0]   io_i_dispatch_packs_1_phy_rs2,
  input  [4:0]   io_i_dispatch_packs_1_arch_rs2,
  input  [6:0]   io_i_dispatch_packs_1_rob_idx,
  input  [63:0]  io_i_dispatch_packs_1_imm,
  input  [63:0]  io_i_dispatch_packs_1_src1_value,
  input  [63:0]  io_i_dispatch_packs_1_src2_value,
  input  [2:0]   io_i_dispatch_packs_1_op1_sel,
  input  [2:0]   io_i_dispatch_packs_1_op2_sel,
  input  [4:0]   io_i_dispatch_packs_1_alu_sel,
  input  [3:0]   io_i_dispatch_packs_1_branch_type,
  input  [1:0]   io_i_dispatch_packs_1_mem_type,
  output         io_o_issue_packs_0_valid,
  output [31:0]  io_o_issue_packs_0_pc,
  output [31:0]  io_o_issue_packs_0_inst,
  output [6:0]   io_o_issue_packs_0_func_code,
  output         io_o_issue_packs_0_branch_predict_pack_valid,
  output [63:0]  io_o_issue_packs_0_branch_predict_pack_target,
  output [3:0]   io_o_issue_packs_0_branch_predict_pack_branch_type,
  output         io_o_issue_packs_0_branch_predict_pack_select,
  output         io_o_issue_packs_0_branch_predict_pack_taken,
  output [6:0]   io_o_issue_packs_0_phy_dst,
  output [6:0]   io_o_issue_packs_0_stale_dst,
  output [4:0]   io_o_issue_packs_0_arch_dst,
  output [2:0]   io_o_issue_packs_0_inst_type,
  output         io_o_issue_packs_0_regWen,
  output         io_o_issue_packs_0_src1_valid,
  output [6:0]   io_o_issue_packs_0_phy_rs1,
  output [4:0]   io_o_issue_packs_0_arch_rs1,
  output         io_o_issue_packs_0_src2_valid,
  output [6:0]   io_o_issue_packs_0_phy_rs2,
  output [4:0]   io_o_issue_packs_0_arch_rs2,
  output [6:0]   io_o_issue_packs_0_rob_idx,
  output [63:0]  io_o_issue_packs_0_imm,
  output [63:0]  io_o_issue_packs_0_src1_value,
  output [63:0]  io_o_issue_packs_0_src2_value,
  output [2:0]   io_o_issue_packs_0_op1_sel,
  output [2:0]   io_o_issue_packs_0_op2_sel,
  output [4:0]   io_o_issue_packs_0_alu_sel,
  output [3:0]   io_o_issue_packs_0_branch_type,
  output [1:0]   io_o_issue_packs_0_mem_type,
  output         io_o_issue_packs_1_valid,
  output [31:0]  io_o_issue_packs_1_pc,
  output [31:0]  io_o_issue_packs_1_inst,
  output [6:0]   io_o_issue_packs_1_func_code,
  output         io_o_issue_packs_1_branch_predict_pack_valid,
  output [63:0]  io_o_issue_packs_1_branch_predict_pack_target,
  output [3:0]   io_o_issue_packs_1_branch_predict_pack_branch_type,
  output         io_o_issue_packs_1_branch_predict_pack_select,
  output         io_o_issue_packs_1_branch_predict_pack_taken,
  output [6:0]   io_o_issue_packs_1_phy_dst,
  output [6:0]   io_o_issue_packs_1_stale_dst,
  output [4:0]   io_o_issue_packs_1_arch_dst,
  output [2:0]   io_o_issue_packs_1_inst_type,
  output         io_o_issue_packs_1_regWen,
  output         io_o_issue_packs_1_src1_valid,
  output [6:0]   io_o_issue_packs_1_phy_rs1,
  output [4:0]   io_o_issue_packs_1_arch_rs1,
  output         io_o_issue_packs_1_src2_valid,
  output [6:0]   io_o_issue_packs_1_phy_rs2,
  output [4:0]   io_o_issue_packs_1_arch_rs2,
  output [6:0]   io_o_issue_packs_1_rob_idx,
  output [63:0]  io_o_issue_packs_1_imm,
  output [63:0]  io_o_issue_packs_1_src1_value,
  output [63:0]  io_o_issue_packs_1_src2_value,
  output [2:0]   io_o_issue_packs_1_op1_sel,
  output [2:0]   io_o_issue_packs_1_op2_sel,
  output [4:0]   io_o_issue_packs_1_alu_sel,
  output [3:0]   io_o_issue_packs_1_branch_type,
  output [1:0]   io_o_issue_packs_1_mem_type,
  input  [127:0] io_i_wakeup_port,
  input          io_i_ex_res_packs_0_valid,
  input  [6:0]   io_i_ex_res_packs_0_uop_func_code,
  input  [6:0]   io_i_ex_res_packs_0_uop_phy_dst,
  input  [63:0]  io_i_ex_res_packs_0_uop_dst_value,
  input          io_i_ex_res_packs_1_valid,
  input  [6:0]   io_i_ex_res_packs_1_uop_func_code,
  input  [6:0]   io_i_ex_res_packs_1_uop_phy_dst,
  input  [63:0]  io_i_ex_res_packs_1_uop_dst_value,
  input          io_i_branch_resolve_pack_valid,
  input          io_i_branch_resolve_pack_mispred,
  input  [6:0]   io_i_branch_resolve_pack_rob_idx,
  output         io_o_full,
  input          io_i_exception,
  input          io_i_rollback_valid,
  input  [1:0]   io_i_available_funcs_0,
  input  [1:0]   io_i_available_funcs_1,
  input  [1:0]   io_i_available_funcs_2,
  input  [1:0]   io_i_available_funcs_3,
  input  [1:0]   io_i_available_funcs_4,
  input  [1:0]   io_i_available_funcs_5,
  input  [6:0]   io_i_ROB_first_entry
);
  wire  reservation_station_0_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_0_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_0_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_0_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_0_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_0_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_0_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_0_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_0_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_0_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_0_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_0_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_0_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_0_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_0_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_0_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_0_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_0_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_0_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_0_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_0_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_0_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_0_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_0_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_0_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_0_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_0_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_0_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_1_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_1_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_1_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_1_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_1_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_1_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_1_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_1_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_1_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_1_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_1_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_1_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_1_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_1_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_1_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_1_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_1_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_1_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_1_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_1_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_1_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_1_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_1_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_1_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_1_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_1_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_1_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_1_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_2_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_2_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_2_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_2_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_2_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_2_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_2_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_2_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_2_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_2_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_2_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_2_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_2_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_2_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_2_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_2_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_2_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_2_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_2_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_2_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_2_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_2_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_2_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_2_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_2_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_2_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_2_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_2_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_3_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_3_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_3_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_3_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_3_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_3_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_3_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_3_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_3_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_3_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_3_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_3_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_3_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_3_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_3_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_3_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_3_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_3_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_3_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_3_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_3_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_3_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_3_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_3_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_3_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_3_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_3_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_3_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_4_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_4_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_4_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_4_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_4_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_4_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_4_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_4_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_4_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_4_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_4_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_4_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_4_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_4_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_4_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_4_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_4_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_4_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_4_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_4_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_4_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_4_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_4_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_4_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_4_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_4_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_4_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_4_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_5_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_5_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_5_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_5_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_5_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_5_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_5_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_5_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_5_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_5_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_5_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_5_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_5_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_5_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_5_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_5_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_5_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_5_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_5_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_5_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_5_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_5_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_5_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_5_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_5_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_5_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_5_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_5_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_6_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_6_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_6_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_6_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_6_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_6_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_6_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_6_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_6_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_6_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_6_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_6_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_6_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_6_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_6_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_6_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_6_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_6_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_6_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_6_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_6_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_6_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_6_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_6_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_6_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_6_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_6_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_6_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_7_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_7_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_7_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_7_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_7_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_7_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_7_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_7_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_7_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_7_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_7_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_7_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_7_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_7_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_7_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_7_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_7_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_7_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_7_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_7_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_7_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_7_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_7_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_7_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_7_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_7_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_7_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_7_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_8_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_8_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_8_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_8_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_8_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_8_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_8_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_8_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_8_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_8_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_8_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_8_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_8_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_8_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_8_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_8_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_8_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_8_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_8_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_8_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_8_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_8_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_8_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_8_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_8_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_8_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_8_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_8_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_9_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_9_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_9_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_9_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_9_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_9_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_9_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_9_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_9_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_9_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_9_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_9_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_9_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_9_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_9_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_9_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_9_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_9_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_9_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_9_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_9_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_9_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_9_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_9_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_9_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_9_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_9_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_9_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_10_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_10_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_10_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_10_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_10_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_10_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_10_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_10_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_10_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_10_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_10_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_10_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_10_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_10_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_10_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_10_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_10_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_10_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_10_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_10_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_10_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_10_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_10_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_10_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_10_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_10_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_10_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_10_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_11_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_11_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_11_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_11_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_11_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_11_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_11_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_11_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_11_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_11_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_11_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_11_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_11_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_11_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_11_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_11_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_11_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_11_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_11_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_11_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_11_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_11_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_11_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_11_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_11_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_11_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_11_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_11_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_12_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_12_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_12_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_12_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_12_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_12_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_12_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_12_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_12_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_12_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_12_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_12_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_12_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_12_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_12_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_12_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_12_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_12_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_12_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_12_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_12_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_12_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_12_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_12_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_12_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_12_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_12_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_12_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_13_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_13_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_13_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_13_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_13_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_13_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_13_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_13_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_13_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_13_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_13_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_13_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_13_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_13_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_13_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_13_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_13_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_13_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_13_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_13_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_13_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_13_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_13_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_13_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_13_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_13_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_13_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_13_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_14_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_14_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_14_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_14_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_14_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_14_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_14_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_14_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_14_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_14_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_14_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_14_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_14_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_14_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_14_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_14_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_14_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_14_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_14_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_14_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_14_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_14_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_14_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_14_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_14_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_14_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_14_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_14_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_15_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_15_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_15_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_15_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_15_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_15_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_15_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_15_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_15_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_15_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_15_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_15_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_15_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_15_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_15_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_15_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_15_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_15_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_15_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_15_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_15_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_15_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_15_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_15_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_15_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_15_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_15_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_15_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_16_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_16_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_16_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_16_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_16_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_16_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_16_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_16_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_16_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_16_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_16_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_16_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_16_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_16_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_16_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_16_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_16_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_16_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_16_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_16_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_16_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_16_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_16_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_16_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_16_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_16_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_16_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_16_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_17_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_17_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_17_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_17_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_17_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_17_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_17_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_17_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_17_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_17_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_17_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_17_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_17_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_17_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_17_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_17_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_17_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_17_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_17_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_17_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_17_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_17_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_17_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_17_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_17_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_17_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_17_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_17_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_18_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_18_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_18_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_18_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_18_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_18_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_18_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_18_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_18_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_18_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_18_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_18_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_18_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_18_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_18_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_18_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_18_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_18_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_18_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_18_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_18_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_18_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_18_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_18_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_18_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_18_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_18_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_18_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_19_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_19_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_19_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_19_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_19_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_19_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_19_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_19_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_19_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_19_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_19_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_19_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_19_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_19_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_19_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_19_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_19_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_19_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_19_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_19_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_19_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_19_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_19_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_19_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_19_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_19_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_19_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_19_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_20_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_20_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_20_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_20_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_20_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_20_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_20_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_20_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_20_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_20_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_20_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_20_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_20_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_20_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_20_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_20_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_20_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_20_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_20_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_20_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_20_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_20_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_20_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_20_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_20_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_20_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_20_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_20_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_21_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_21_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_21_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_21_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_21_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_21_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_21_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_21_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_21_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_21_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_21_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_21_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_21_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_21_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_21_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_21_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_21_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_21_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_21_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_21_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_21_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_21_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_21_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_21_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_21_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_21_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_21_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_21_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_22_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_22_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_22_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_22_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_22_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_22_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_22_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_22_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_22_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_22_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_22_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_22_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_22_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_22_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_22_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_22_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_22_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_22_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_22_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_22_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_22_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_22_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_22_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_22_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_22_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_22_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_22_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_22_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_23_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_23_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_23_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_23_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_23_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_23_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_23_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_23_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_23_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_23_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_23_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_23_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_23_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_23_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_23_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_23_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_23_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_23_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_23_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_23_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_23_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_23_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_23_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_23_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_23_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_23_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_23_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_23_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_24_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_24_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_24_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_24_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_24_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_24_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_24_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_24_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_24_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_24_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_24_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_24_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_24_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_24_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_24_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_24_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_24_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_24_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_24_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_24_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_24_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_24_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_24_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_24_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_24_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_24_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_24_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_24_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_25_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_25_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_25_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_25_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_25_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_25_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_25_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_25_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_25_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_25_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_25_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_25_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_25_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_25_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_25_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_25_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_25_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_25_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_25_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_25_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_25_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_25_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_25_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_25_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_25_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_25_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_25_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_25_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_26_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_26_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_26_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_26_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_26_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_26_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_26_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_26_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_26_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_26_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_26_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_26_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_26_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_26_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_26_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_26_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_26_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_26_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_26_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_26_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_26_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_26_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_26_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_26_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_26_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_26_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_26_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_26_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_27_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_27_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_27_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_27_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_27_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_27_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_27_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_27_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_27_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_27_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_27_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_27_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_27_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_27_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_27_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_27_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_27_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_27_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_27_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_27_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_27_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_27_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_27_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_27_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_27_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_27_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_27_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_27_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_28_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_28_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_28_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_28_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_28_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_28_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_28_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_28_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_28_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_28_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_28_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_28_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_28_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_28_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_28_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_28_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_28_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_28_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_28_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_28_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_28_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_28_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_28_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_28_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_28_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_28_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_28_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_28_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_29_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_29_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_29_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_29_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_29_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_29_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_29_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_29_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_29_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_29_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_29_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_29_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_29_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_29_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_29_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_29_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_29_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_29_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_29_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_29_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_29_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_29_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_29_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_29_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_29_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_29_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_29_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_29_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_30_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_30_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_30_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_30_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_30_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_30_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_30_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_30_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_30_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_30_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_30_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_30_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_30_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_30_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_30_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_30_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_30_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_30_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_30_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_30_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_30_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_30_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_30_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_30_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_30_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_30_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_30_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_30_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_clock; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_reset; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_o_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_o_ready_to_issue; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_issue_granted; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_exception; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_write_slot; // @[reservation_station.scala 38:56]
  wire [127:0] reservation_station_31_io_i_wakeup_port; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_uop_valid; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_31_io_i_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_31_io_i_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_31_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_31_io_i_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_31_io_i_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_31_io_i_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_i_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_31_io_i_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_i_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_i_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_i_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_31_io_i_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_31_io_i_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_31_io_i_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_31_io_i_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_31_io_i_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_31_io_o_uop_pc; // @[reservation_station.scala 38:56]
  wire [31:0] reservation_station_31_io_o_uop_inst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_o_uop_func_code; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_31_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_o_uop_phy_dst; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_o_uop_stale_dst; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_31_io_o_uop_arch_dst; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_31_io_o_uop_inst_type; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_o_uop_regWen; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_o_uop_src1_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_o_uop_phy_rs1; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_31_io_o_uop_arch_rs1; // @[reservation_station.scala 38:56]
  wire  reservation_station_31_io_o_uop_src2_valid; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_o_uop_phy_rs2; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_31_io_o_uop_arch_rs2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_o_uop_rob_idx; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_o_uop_imm; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_o_uop_src1_value; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_o_uop_src2_value; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_31_io_o_uop_op1_sel; // @[reservation_station.scala 38:56]
  wire [2:0] reservation_station_31_io_o_uop_op2_sel; // @[reservation_station.scala 38:56]
  wire [4:0] reservation_station_31_io_o_uop_alu_sel; // @[reservation_station.scala 38:56]
  wire [3:0] reservation_station_31_io_o_uop_branch_type; // @[reservation_station.scala 38:56]
  wire [1:0] reservation_station_31_io_o_uop_mem_type; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_exe_dst1; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_exe_dst2; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_i_exe_value1; // @[reservation_station.scala 38:56]
  wire [63:0] reservation_station_31_io_i_exe_value2; // @[reservation_station.scala 38:56]
  wire [6:0] reservation_station_31_io_i_ROB_first_entry; // @[reservation_station.scala 38:56]
  wire  temp_1 = reservation_station_1_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_0 = reservation_station_0_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_3 = reservation_station_3_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_2 = reservation_station_2_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_5 = reservation_station_5_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_4 = reservation_station_4_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_7 = reservation_station_7_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_6 = reservation_station_6_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_lo_lo = {temp_7,temp_6,temp_5,temp_4,temp_3,temp_2,temp_1,temp_0}; // @[reservation_station.scala 48:46]
  wire  temp_9 = reservation_station_9_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_8 = reservation_station_8_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_11 = reservation_station_11_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_10 = reservation_station_10_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_13 = reservation_station_13_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_12 = reservation_station_12_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_15 = reservation_station_15_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_14 = reservation_station_14_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [15:0] reservation_station_valid_lo = {temp_15,temp_14,temp_13,temp_12,temp_11,temp_10,temp_9,temp_8,
    reservation_station_valid_lo_lo}; // @[reservation_station.scala 48:46]
  wire  temp_17 = reservation_station_17_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_16 = reservation_station_16_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_19 = reservation_station_19_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_18 = reservation_station_18_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_21 = reservation_station_21_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_20 = reservation_station_20_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_23 = reservation_station_23_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_22 = reservation_station_22_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_hi_lo = {temp_23,temp_22,temp_21,temp_20,temp_19,temp_18,temp_17,temp_16}; // @[reservation_station.scala 48:46]
  wire  temp_25 = reservation_station_25_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_24 = reservation_station_24_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_27 = reservation_station_27_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_26 = reservation_station_26_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_29 = reservation_station_29_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_28 = reservation_station_28_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_31 = reservation_station_31_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_30 = reservation_station_30_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [31:0] reservation_station_valid = {temp_31,temp_30,temp_29,temp_28,temp_27,temp_26,temp_25,temp_24,
    reservation_station_valid_hi_lo,reservation_station_valid_lo}; // @[reservation_station.scala 48:46]
  wire [31:0] _write_idx1_T = ~reservation_station_valid; // @[reservation_station.scala 49:34]
  wire [4:0] _write_idx1_T_33 = _write_idx1_T[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_34 = _write_idx1_T[29] ? 5'h1d : _write_idx1_T_33; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_35 = _write_idx1_T[28] ? 5'h1c : _write_idx1_T_34; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_36 = _write_idx1_T[27] ? 5'h1b : _write_idx1_T_35; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_37 = _write_idx1_T[26] ? 5'h1a : _write_idx1_T_36; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_38 = _write_idx1_T[25] ? 5'h19 : _write_idx1_T_37; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_39 = _write_idx1_T[24] ? 5'h18 : _write_idx1_T_38; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_40 = _write_idx1_T[23] ? 5'h17 : _write_idx1_T_39; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_41 = _write_idx1_T[22] ? 5'h16 : _write_idx1_T_40; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_42 = _write_idx1_T[21] ? 5'h15 : _write_idx1_T_41; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_43 = _write_idx1_T[20] ? 5'h14 : _write_idx1_T_42; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_44 = _write_idx1_T[19] ? 5'h13 : _write_idx1_T_43; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_45 = _write_idx1_T[18] ? 5'h12 : _write_idx1_T_44; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_46 = _write_idx1_T[17] ? 5'h11 : _write_idx1_T_45; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_47 = _write_idx1_T[16] ? 5'h10 : _write_idx1_T_46; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_48 = _write_idx1_T[15] ? 5'hf : _write_idx1_T_47; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_49 = _write_idx1_T[14] ? 5'he : _write_idx1_T_48; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_50 = _write_idx1_T[13] ? 5'hd : _write_idx1_T_49; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_51 = _write_idx1_T[12] ? 5'hc : _write_idx1_T_50; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_52 = _write_idx1_T[11] ? 5'hb : _write_idx1_T_51; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_53 = _write_idx1_T[10] ? 5'ha : _write_idx1_T_52; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_54 = _write_idx1_T[9] ? 5'h9 : _write_idx1_T_53; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_55 = _write_idx1_T[8] ? 5'h8 : _write_idx1_T_54; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_56 = _write_idx1_T[7] ? 5'h7 : _write_idx1_T_55; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_57 = _write_idx1_T[6] ? 5'h6 : _write_idx1_T_56; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_58 = _write_idx1_T[5] ? 5'h5 : _write_idx1_T_57; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_59 = _write_idx1_T[4] ? 5'h4 : _write_idx1_T_58; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_60 = _write_idx1_T[3] ? 5'h3 : _write_idx1_T_59; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_61 = _write_idx1_T[2] ? 5'h2 : _write_idx1_T_60; // @[Mux.scala 47:70]
  wire [4:0] _write_idx1_T_62 = _write_idx1_T[1] ? 5'h1 : _write_idx1_T_61; // @[Mux.scala 47:70]
  wire [4:0] write_idx1 = _write_idx1_T[0] ? 5'h0 : _write_idx1_T_62; // @[Mux.scala 47:70]
  wire [31:0] _reservation_station_valid_withmask_T = 32'h1 << write_idx1; // @[OneHot.scala 57:35]
  wire [31:0] reservation_station_valid_withmask = reservation_station_valid | _reservation_station_valid_withmask_T; // @[reservation_station.scala 50:69]
  wire [31:0] _write_idx2_T = ~reservation_station_valid_withmask; // @[reservation_station.scala 51:34]
  wire [4:0] _write_idx2_T_33 = _write_idx2_T[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_34 = _write_idx2_T[29] ? 5'h1d : _write_idx2_T_33; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_35 = _write_idx2_T[28] ? 5'h1c : _write_idx2_T_34; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_36 = _write_idx2_T[27] ? 5'h1b : _write_idx2_T_35; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_37 = _write_idx2_T[26] ? 5'h1a : _write_idx2_T_36; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_38 = _write_idx2_T[25] ? 5'h19 : _write_idx2_T_37; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_39 = _write_idx2_T[24] ? 5'h18 : _write_idx2_T_38; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_40 = _write_idx2_T[23] ? 5'h17 : _write_idx2_T_39; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_41 = _write_idx2_T[22] ? 5'h16 : _write_idx2_T_40; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_42 = _write_idx2_T[21] ? 5'h15 : _write_idx2_T_41; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_43 = _write_idx2_T[20] ? 5'h14 : _write_idx2_T_42; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_44 = _write_idx2_T[19] ? 5'h13 : _write_idx2_T_43; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_45 = _write_idx2_T[18] ? 5'h12 : _write_idx2_T_44; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_46 = _write_idx2_T[17] ? 5'h11 : _write_idx2_T_45; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_47 = _write_idx2_T[16] ? 5'h10 : _write_idx2_T_46; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_48 = _write_idx2_T[15] ? 5'hf : _write_idx2_T_47; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_49 = _write_idx2_T[14] ? 5'he : _write_idx2_T_48; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_50 = _write_idx2_T[13] ? 5'hd : _write_idx2_T_49; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_51 = _write_idx2_T[12] ? 5'hc : _write_idx2_T_50; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_52 = _write_idx2_T[11] ? 5'hb : _write_idx2_T_51; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_53 = _write_idx2_T[10] ? 5'ha : _write_idx2_T_52; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_54 = _write_idx2_T[9] ? 5'h9 : _write_idx2_T_53; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_55 = _write_idx2_T[8] ? 5'h8 : _write_idx2_T_54; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_56 = _write_idx2_T[7] ? 5'h7 : _write_idx2_T_55; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_57 = _write_idx2_T[6] ? 5'h6 : _write_idx2_T_56; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_58 = _write_idx2_T[5] ? 5'h5 : _write_idx2_T_57; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_59 = _write_idx2_T[4] ? 5'h4 : _write_idx2_T_58; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_60 = _write_idx2_T[3] ? 5'h3 : _write_idx2_T_59; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_61 = _write_idx2_T[2] ? 5'h2 : _write_idx2_T_60; // @[Mux.scala 47:70]
  wire [4:0] _write_idx2_T_62 = _write_idx2_T[1] ? 5'h1 : _write_idx2_T_61; // @[Mux.scala 47:70]
  wire [4:0] write_idx2 = _write_idx2_T[0] ? 5'h0 : _write_idx2_T_62; // @[Mux.scala 47:70]
  wire  temp2_0 = |io_i_available_funcs_0; // @[reservation_station.scala 59:44]
  wire  temp2_1 = |io_i_available_funcs_1; // @[reservation_station.scala 59:44]
  wire  temp2_2 = |io_i_available_funcs_2; // @[reservation_station.scala 59:44]
  wire  temp2_3 = |io_i_available_funcs_3; // @[reservation_station.scala 59:44]
  wire  temp2_4 = |io_i_available_funcs_4; // @[reservation_station.scala 59:44]
  wire  temp2_5 = |io_i_available_funcs_5; // @[reservation_station.scala 59:44]
  wire [6:0] available_funcs = {1'h0,temp2_5,temp2_4,temp2_3,temp2_2,temp2_1,temp2_0}; // @[reservation_station.scala 61:37]
  wire [6:0] _slots_can_issue_T = reservation_station_0_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_0 = reservation_station_0_io_o_ready_to_issue & |_slots_can_issue_T; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_4 = reservation_station_1_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_1 = reservation_station_1_io_o_ready_to_issue & |_slots_can_issue_T_4; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_8 = reservation_station_2_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_2 = reservation_station_2_io_o_ready_to_issue & |_slots_can_issue_T_8; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_12 = reservation_station_3_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_3 = reservation_station_3_io_o_ready_to_issue & |_slots_can_issue_T_12; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_16 = reservation_station_4_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_4 = reservation_station_4_io_o_ready_to_issue & |_slots_can_issue_T_16; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_20 = reservation_station_5_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_5 = reservation_station_5_io_o_ready_to_issue & |_slots_can_issue_T_20; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_24 = reservation_station_6_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_6 = reservation_station_6_io_o_ready_to_issue & |_slots_can_issue_T_24; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_28 = reservation_station_7_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_7 = reservation_station_7_io_o_ready_to_issue & |_slots_can_issue_T_28; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_32 = reservation_station_8_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_8 = reservation_station_8_io_o_ready_to_issue & |_slots_can_issue_T_32; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_36 = reservation_station_9_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_9 = reservation_station_9_io_o_ready_to_issue & |_slots_can_issue_T_36; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_40 = reservation_station_10_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_10 = reservation_station_10_io_o_ready_to_issue & |_slots_can_issue_T_40; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_44 = reservation_station_11_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_11 = reservation_station_11_io_o_ready_to_issue & |_slots_can_issue_T_44; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_48 = reservation_station_12_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_12 = reservation_station_12_io_o_ready_to_issue & |_slots_can_issue_T_48; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_52 = reservation_station_13_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_13 = reservation_station_13_io_o_ready_to_issue & |_slots_can_issue_T_52; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_56 = reservation_station_14_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_14 = reservation_station_14_io_o_ready_to_issue & |_slots_can_issue_T_56; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_60 = reservation_station_15_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_15 = reservation_station_15_io_o_ready_to_issue & |_slots_can_issue_T_60; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_64 = reservation_station_16_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_16 = reservation_station_16_io_o_ready_to_issue & |_slots_can_issue_T_64; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_68 = reservation_station_17_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_17 = reservation_station_17_io_o_ready_to_issue & |_slots_can_issue_T_68; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_72 = reservation_station_18_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_18 = reservation_station_18_io_o_ready_to_issue & |_slots_can_issue_T_72; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_76 = reservation_station_19_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_19 = reservation_station_19_io_o_ready_to_issue & |_slots_can_issue_T_76; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_80 = reservation_station_20_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_20 = reservation_station_20_io_o_ready_to_issue & |_slots_can_issue_T_80; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_84 = reservation_station_21_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_21 = reservation_station_21_io_o_ready_to_issue & |_slots_can_issue_T_84; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_88 = reservation_station_22_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_22 = reservation_station_22_io_o_ready_to_issue & |_slots_can_issue_T_88; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_92 = reservation_station_23_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_23 = reservation_station_23_io_o_ready_to_issue & |_slots_can_issue_T_92; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_96 = reservation_station_24_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_24 = reservation_station_24_io_o_ready_to_issue & |_slots_can_issue_T_96; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_100 = reservation_station_25_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_25 = reservation_station_25_io_o_ready_to_issue & |_slots_can_issue_T_100; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_104 = reservation_station_26_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_26 = reservation_station_26_io_o_ready_to_issue & |_slots_can_issue_T_104; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_108 = reservation_station_27_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_27 = reservation_station_27_io_o_ready_to_issue & |_slots_can_issue_T_108; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_112 = reservation_station_28_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_28 = reservation_station_28_io_o_ready_to_issue & |_slots_can_issue_T_112; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_116 = reservation_station_29_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_29 = reservation_station_29_io_o_ready_to_issue & |_slots_can_issue_T_116; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_120 = reservation_station_30_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_30 = reservation_station_30_io_o_ready_to_issue & |_slots_can_issue_T_120; // @[reservation_station.scala 63:103]
  wire [6:0] _slots_can_issue_T_124 = reservation_station_31_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:150]
  wire  slots_can_issue_31 = reservation_station_31_io_o_ready_to_issue & |_slots_can_issue_T_124; // @[reservation_station.scala 63:103]
  wire [7:0] issue1_idx_lo_lo = {slots_can_issue_7,slots_can_issue_6,slots_can_issue_5,slots_can_issue_4,
    slots_can_issue_3,slots_can_issue_2,slots_can_issue_1,slots_can_issue_0}; // @[reservation_station.scala 65:58]
  wire [15:0] issue1_idx_lo = {slots_can_issue_15,slots_can_issue_14,slots_can_issue_13,slots_can_issue_12,
    slots_can_issue_11,slots_can_issue_10,slots_can_issue_9,slots_can_issue_8,issue1_idx_lo_lo}; // @[reservation_station.scala 65:58]
  wire [7:0] issue1_idx_hi_lo = {slots_can_issue_23,slots_can_issue_22,slots_can_issue_21,slots_can_issue_20,
    slots_can_issue_19,slots_can_issue_18,slots_can_issue_17,slots_can_issue_16}; // @[reservation_station.scala 65:58]
  wire [31:0] _issue1_idx_T = {slots_can_issue_31,slots_can_issue_30,slots_can_issue_29,slots_can_issue_28,
    slots_can_issue_27,slots_can_issue_26,slots_can_issue_25,slots_can_issue_24,issue1_idx_hi_lo,issue1_idx_lo}; // @[reservation_station.scala 65:58]
  wire [4:0] _issue1_idx_T_33 = _issue1_idx_T[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_34 = _issue1_idx_T[29] ? 5'h1d : _issue1_idx_T_33; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_35 = _issue1_idx_T[28] ? 5'h1c : _issue1_idx_T_34; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_36 = _issue1_idx_T[27] ? 5'h1b : _issue1_idx_T_35; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_37 = _issue1_idx_T[26] ? 5'h1a : _issue1_idx_T_36; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_38 = _issue1_idx_T[25] ? 5'h19 : _issue1_idx_T_37; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_39 = _issue1_idx_T[24] ? 5'h18 : _issue1_idx_T_38; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_40 = _issue1_idx_T[23] ? 5'h17 : _issue1_idx_T_39; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_41 = _issue1_idx_T[22] ? 5'h16 : _issue1_idx_T_40; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_42 = _issue1_idx_T[21] ? 5'h15 : _issue1_idx_T_41; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_43 = _issue1_idx_T[20] ? 5'h14 : _issue1_idx_T_42; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_44 = _issue1_idx_T[19] ? 5'h13 : _issue1_idx_T_43; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_45 = _issue1_idx_T[18] ? 5'h12 : _issue1_idx_T_44; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_46 = _issue1_idx_T[17] ? 5'h11 : _issue1_idx_T_45; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_47 = _issue1_idx_T[16] ? 5'h10 : _issue1_idx_T_46; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_48 = _issue1_idx_T[15] ? 5'hf : _issue1_idx_T_47; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_49 = _issue1_idx_T[14] ? 5'he : _issue1_idx_T_48; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_50 = _issue1_idx_T[13] ? 5'hd : _issue1_idx_T_49; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_51 = _issue1_idx_T[12] ? 5'hc : _issue1_idx_T_50; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_52 = _issue1_idx_T[11] ? 5'hb : _issue1_idx_T_51; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_53 = _issue1_idx_T[10] ? 5'ha : _issue1_idx_T_52; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_54 = _issue1_idx_T[9] ? 5'h9 : _issue1_idx_T_53; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_55 = _issue1_idx_T[8] ? 5'h8 : _issue1_idx_T_54; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_56 = _issue1_idx_T[7] ? 5'h7 : _issue1_idx_T_55; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_57 = _issue1_idx_T[6] ? 5'h6 : _issue1_idx_T_56; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_58 = _issue1_idx_T[5] ? 5'h5 : _issue1_idx_T_57; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_59 = _issue1_idx_T[4] ? 5'h4 : _issue1_idx_T_58; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_60 = _issue1_idx_T[3] ? 5'h3 : _issue1_idx_T_59; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_61 = _issue1_idx_T[2] ? 5'h2 : _issue1_idx_T_60; // @[Mux.scala 47:70]
  wire [4:0] _issue1_idx_T_62 = _issue1_idx_T[1] ? 5'h1 : _issue1_idx_T_61; // @[Mux.scala 47:70]
  wire [4:0] issue1_idx = _issue1_idx_T[0] ? 5'h0 : _issue1_idx_T_62; // @[Mux.scala 47:70]
  wire  _issue1_func_code_T = 5'h0 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_1 = 5'h1 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_2 = 5'h2 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_3 = 5'h3 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_4 = 5'h4 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_5 = 5'h5 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_6 = 5'h6 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_7 = 5'h7 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_8 = 5'h8 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_9 = 5'h9 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_10 = 5'ha == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_11 = 5'hb == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_12 = 5'hc == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_13 = 5'hd == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_14 = 5'he == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_15 = 5'hf == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_16 = 5'h10 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_17 = 5'h11 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_18 = 5'h12 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_19 = 5'h13 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_20 = 5'h14 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_21 = 5'h15 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_22 = 5'h16 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_23 = 5'h17 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_24 = 5'h18 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_25 = 5'h19 == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_26 = 5'h1a == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_27 = 5'h1b == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_28 = 5'h1c == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_29 = 5'h1d == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_30 = 5'h1e == issue1_idx; // @[reservation_station.scala 68:85]
  wire  _issue1_func_code_T_31 = 5'h1f == issue1_idx; // @[reservation_station.scala 68:85]
  wire [6:0] _issue1_func_code_T_32 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_func_code : 7'h40; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_33 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_func_code :
    _issue1_func_code_T_32; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_34 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_func_code :
    _issue1_func_code_T_33; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_35 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_func_code :
    _issue1_func_code_T_34; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_36 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_func_code :
    _issue1_func_code_T_35; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_37 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_func_code :
    _issue1_func_code_T_36; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_38 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_func_code :
    _issue1_func_code_T_37; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_39 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_func_code :
    _issue1_func_code_T_38; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_40 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_func_code :
    _issue1_func_code_T_39; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_41 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_func_code :
    _issue1_func_code_T_40; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_42 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_func_code :
    _issue1_func_code_T_41; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_43 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_func_code :
    _issue1_func_code_T_42; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_44 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_func_code :
    _issue1_func_code_T_43; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_45 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_func_code :
    _issue1_func_code_T_44; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_46 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_func_code :
    _issue1_func_code_T_45; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_47 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_func_code :
    _issue1_func_code_T_46; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_48 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_func_code :
    _issue1_func_code_T_47; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_49 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_func_code :
    _issue1_func_code_T_48; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_50 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_func_code :
    _issue1_func_code_T_49; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_51 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_func_code :
    _issue1_func_code_T_50; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_52 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_func_code :
    _issue1_func_code_T_51; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_53 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_func_code :
    _issue1_func_code_T_52; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_54 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_func_code :
    _issue1_func_code_T_53; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_55 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_func_code :
    _issue1_func_code_T_54; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_56 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_func_code :
    _issue1_func_code_T_55; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_57 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_func_code :
    _issue1_func_code_T_56; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_58 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_func_code :
    _issue1_func_code_T_57; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_59 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_func_code :
    _issue1_func_code_T_58; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_60 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_func_code :
    _issue1_func_code_T_59; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_61 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_func_code :
    _issue1_func_code_T_60; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_62 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_func_code :
    _issue1_func_code_T_61; // @[Mux.scala 101:16]
  wire [6:0] issue1_func_code = _issue1_func_code_T ? reservation_station_0_io_o_uop_func_code : _issue1_func_code_T_62; // @[Mux.scala 101:16]
  wire [2:0] hi = issue1_func_code[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] lo = issue1_func_code[3:0]; // @[OneHot.scala 31:18]
  wire  _T = |hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_14 = {{1'd0}, hi}; // @[OneHot.scala 32:28]
  wire [3:0] _T_1 = _GEN_14 | lo; // @[OneHot.scala 32:28]
  wire [1:0] hi_1 = _T_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_1 = _T_1[1:0]; // @[OneHot.scala 31:18]
  wire  _T_2 = |hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _T_3 = hi_1 | lo_1; // @[OneHot.scala 32:28]
  wire [2:0] _T_6 = {_T,_T_2,_T_3[1]}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_1 = 3'h1 == _T_6 ? io_i_available_funcs_1 : io_i_available_funcs_0; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_2 = 3'h2 == _T_6 ? io_i_available_funcs_2 : _GEN_1; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_3 = 3'h3 == _T_6 ? io_i_available_funcs_3 : _GEN_2; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_4 = 3'h4 == _T_6 ? io_i_available_funcs_4 : _GEN_3; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_5 = 3'h5 == _T_6 ? io_i_available_funcs_5 : _GEN_4; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_6 = 3'h6 == _T_6 ? 2'h0 : _GEN_5; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _available_funcs_with_mask_T_8 = _GEN_6 - 2'h1; // @[reservation_station.scala 71:109]
  wire [1:0] available_funcs_with_mask_0 = 3'h0 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_0; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_1 = 3'h1 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_1; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_2 = 3'h2 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_2; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_3 = 3'h3 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_3; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_4 = 3'h4 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_4; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_5 = 3'h5 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_5; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_6 = 3'h6 == _T_6 ? _available_funcs_with_mask_T_8 : 2'h0; // @[reservation_station.scala 70:31 71:{59,59}]
  wire  temp3_0 = |available_funcs_with_mask_0; // @[reservation_station.scala 75:49]
  wire  temp3_1 = |available_funcs_with_mask_1; // @[reservation_station.scala 75:49]
  wire  temp3_2 = |available_funcs_with_mask_2; // @[reservation_station.scala 75:49]
  wire  temp3_3 = |available_funcs_with_mask_3; // @[reservation_station.scala 75:49]
  wire  temp3_4 = |available_funcs_with_mask_4; // @[reservation_station.scala 75:49]
  wire  temp3_5 = |available_funcs_with_mask_5; // @[reservation_station.scala 75:49]
  wire  temp3_6 = |available_funcs_with_mask_6; // @[reservation_station.scala 75:49]
  wire [6:0] available_funcs2_bits = {temp3_6,temp3_5,temp3_4,temp3_3,temp3_2,temp3_1,temp3_0}; // @[reservation_station.scala 78:46]
  wire [6:0] _slots_can_issue2_T_2 = reservation_station_0_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_3 = |_slots_can_issue2_T_2; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_0 = slots_can_issue_0 & 5'h0 != issue1_idx & _slots_can_issue2_T_3; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_8 = reservation_station_1_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_9 = |_slots_can_issue2_T_8; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_1 = slots_can_issue_1 & 5'h1 != issue1_idx & _slots_can_issue2_T_9; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_14 = reservation_station_2_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_15 = |_slots_can_issue2_T_14; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_2 = slots_can_issue_2 & 5'h2 != issue1_idx & _slots_can_issue2_T_15; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_20 = reservation_station_3_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_21 = |_slots_can_issue2_T_20; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_3 = slots_can_issue_3 & 5'h3 != issue1_idx & _slots_can_issue2_T_21; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_26 = reservation_station_4_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_27 = |_slots_can_issue2_T_26; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_4 = slots_can_issue_4 & 5'h4 != issue1_idx & _slots_can_issue2_T_27; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_32 = reservation_station_5_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_33 = |_slots_can_issue2_T_32; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_5 = slots_can_issue_5 & 5'h5 != issue1_idx & _slots_can_issue2_T_33; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_38 = reservation_station_6_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_39 = |_slots_can_issue2_T_38; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_6 = slots_can_issue_6 & 5'h6 != issue1_idx & _slots_can_issue2_T_39; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_44 = reservation_station_7_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_45 = |_slots_can_issue2_T_44; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_7 = slots_can_issue_7 & 5'h7 != issue1_idx & _slots_can_issue2_T_45; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_50 = reservation_station_8_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_51 = |_slots_can_issue2_T_50; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_8 = slots_can_issue_8 & 5'h8 != issue1_idx & _slots_can_issue2_T_51; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_56 = reservation_station_9_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_57 = |_slots_can_issue2_T_56; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_9 = slots_can_issue_9 & 5'h9 != issue1_idx & _slots_can_issue2_T_57; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_62 = reservation_station_10_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_63 = |_slots_can_issue2_T_62; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_10 = slots_can_issue_10 & 5'ha != issue1_idx & _slots_can_issue2_T_63; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_68 = reservation_station_11_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_69 = |_slots_can_issue2_T_68; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_11 = slots_can_issue_11 & 5'hb != issue1_idx & _slots_can_issue2_T_69; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_74 = reservation_station_12_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_75 = |_slots_can_issue2_T_74; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_12 = slots_can_issue_12 & 5'hc != issue1_idx & _slots_can_issue2_T_75; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_80 = reservation_station_13_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_81 = |_slots_can_issue2_T_80; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_13 = slots_can_issue_13 & 5'hd != issue1_idx & _slots_can_issue2_T_81; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_86 = reservation_station_14_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_87 = |_slots_can_issue2_T_86; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_14 = slots_can_issue_14 & 5'he != issue1_idx & _slots_can_issue2_T_87; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_92 = reservation_station_15_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_93 = |_slots_can_issue2_T_92; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_15 = slots_can_issue_15 & 5'hf != issue1_idx & _slots_can_issue2_T_93; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_98 = reservation_station_16_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_99 = |_slots_can_issue2_T_98; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_16 = slots_can_issue_16 & 5'h10 != issue1_idx & _slots_can_issue2_T_99; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_104 = reservation_station_17_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_105 = |_slots_can_issue2_T_104; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_17 = slots_can_issue_17 & 5'h11 != issue1_idx & _slots_can_issue2_T_105; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_110 = reservation_station_18_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_111 = |_slots_can_issue2_T_110; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_18 = slots_can_issue_18 & 5'h12 != issue1_idx & _slots_can_issue2_T_111; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_116 = reservation_station_19_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_117 = |_slots_can_issue2_T_116; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_19 = slots_can_issue_19 & 5'h13 != issue1_idx & _slots_can_issue2_T_117; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_122 = reservation_station_20_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_123 = |_slots_can_issue2_T_122; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_20 = slots_can_issue_20 & 5'h14 != issue1_idx & _slots_can_issue2_T_123; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_128 = reservation_station_21_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_129 = |_slots_can_issue2_T_128; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_21 = slots_can_issue_21 & 5'h15 != issue1_idx & _slots_can_issue2_T_129; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_134 = reservation_station_22_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_135 = |_slots_can_issue2_T_134; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_22 = slots_can_issue_22 & 5'h16 != issue1_idx & _slots_can_issue2_T_135; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_140 = reservation_station_23_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_141 = |_slots_can_issue2_T_140; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_23 = slots_can_issue_23 & 5'h17 != issue1_idx & _slots_can_issue2_T_141; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_146 = reservation_station_24_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_147 = |_slots_can_issue2_T_146; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_24 = slots_can_issue_24 & 5'h18 != issue1_idx & _slots_can_issue2_T_147; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_152 = reservation_station_25_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_153 = |_slots_can_issue2_T_152; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_25 = slots_can_issue_25 & 5'h19 != issue1_idx & _slots_can_issue2_T_153; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_158 = reservation_station_26_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_159 = |_slots_can_issue2_T_158; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_26 = slots_can_issue_26 & 5'h1a != issue1_idx & _slots_can_issue2_T_159; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_164 = reservation_station_27_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_165 = |_slots_can_issue2_T_164; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_27 = slots_can_issue_27 & 5'h1b != issue1_idx & _slots_can_issue2_T_165; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_170 = reservation_station_28_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_171 = |_slots_can_issue2_T_170; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_28 = slots_can_issue_28 & 5'h1c != issue1_idx & _slots_can_issue2_T_171; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_176 = reservation_station_29_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_177 = |_slots_can_issue2_T_176; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_29 = slots_can_issue_29 & 5'h1d != issue1_idx & _slots_can_issue2_T_177; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_182 = reservation_station_30_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_183 = |_slots_can_issue2_T_182; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_30 = slots_can_issue_30 & 5'h1e != issue1_idx & _slots_can_issue2_T_183; // @[reservation_station.scala 79:104]
  wire [6:0] _slots_can_issue2_T_188 = reservation_station_31_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_189 = |_slots_can_issue2_T_188; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_31 = slots_can_issue_31 & 5'h1f != issue1_idx & _slots_can_issue2_T_189; // @[reservation_station.scala 79:104]
  wire [7:0] issue2_idx_lo_lo = {slots_can_issue2_7,slots_can_issue2_6,slots_can_issue2_5,slots_can_issue2_4,
    slots_can_issue2_3,slots_can_issue2_2,slots_can_issue2_1,slots_can_issue2_0}; // @[reservation_station.scala 83:53]
  wire [15:0] issue2_idx_lo = {slots_can_issue2_15,slots_can_issue2_14,slots_can_issue2_13,slots_can_issue2_12,
    slots_can_issue2_11,slots_can_issue2_10,slots_can_issue2_9,slots_can_issue2_8,issue2_idx_lo_lo}; // @[reservation_station.scala 83:53]
  wire [7:0] issue2_idx_hi_lo = {slots_can_issue2_23,slots_can_issue2_22,slots_can_issue2_21,slots_can_issue2_20,
    slots_can_issue2_19,slots_can_issue2_18,slots_can_issue2_17,slots_can_issue2_16}; // @[reservation_station.scala 83:53]
  wire [31:0] _issue2_idx_T = {slots_can_issue2_31,slots_can_issue2_30,slots_can_issue2_29,slots_can_issue2_28,
    slots_can_issue2_27,slots_can_issue2_26,slots_can_issue2_25,slots_can_issue2_24,issue2_idx_hi_lo,issue2_idx_lo}; // @[reservation_station.scala 83:53]
  wire [4:0] _issue2_idx_T_33 = _issue2_idx_T[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_34 = _issue2_idx_T[29] ? 5'h1d : _issue2_idx_T_33; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_35 = _issue2_idx_T[28] ? 5'h1c : _issue2_idx_T_34; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_36 = _issue2_idx_T[27] ? 5'h1b : _issue2_idx_T_35; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_37 = _issue2_idx_T[26] ? 5'h1a : _issue2_idx_T_36; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_38 = _issue2_idx_T[25] ? 5'h19 : _issue2_idx_T_37; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_39 = _issue2_idx_T[24] ? 5'h18 : _issue2_idx_T_38; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_40 = _issue2_idx_T[23] ? 5'h17 : _issue2_idx_T_39; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_41 = _issue2_idx_T[22] ? 5'h16 : _issue2_idx_T_40; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_42 = _issue2_idx_T[21] ? 5'h15 : _issue2_idx_T_41; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_43 = _issue2_idx_T[20] ? 5'h14 : _issue2_idx_T_42; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_44 = _issue2_idx_T[19] ? 5'h13 : _issue2_idx_T_43; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_45 = _issue2_idx_T[18] ? 5'h12 : _issue2_idx_T_44; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_46 = _issue2_idx_T[17] ? 5'h11 : _issue2_idx_T_45; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_47 = _issue2_idx_T[16] ? 5'h10 : _issue2_idx_T_46; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_48 = _issue2_idx_T[15] ? 5'hf : _issue2_idx_T_47; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_49 = _issue2_idx_T[14] ? 5'he : _issue2_idx_T_48; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_50 = _issue2_idx_T[13] ? 5'hd : _issue2_idx_T_49; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_51 = _issue2_idx_T[12] ? 5'hc : _issue2_idx_T_50; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_52 = _issue2_idx_T[11] ? 5'hb : _issue2_idx_T_51; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_53 = _issue2_idx_T[10] ? 5'ha : _issue2_idx_T_52; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_54 = _issue2_idx_T[9] ? 5'h9 : _issue2_idx_T_53; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_55 = _issue2_idx_T[8] ? 5'h8 : _issue2_idx_T_54; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_56 = _issue2_idx_T[7] ? 5'h7 : _issue2_idx_T_55; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_57 = _issue2_idx_T[6] ? 5'h6 : _issue2_idx_T_56; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_58 = _issue2_idx_T[5] ? 5'h5 : _issue2_idx_T_57; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_59 = _issue2_idx_T[4] ? 5'h4 : _issue2_idx_T_58; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_60 = _issue2_idx_T[3] ? 5'h3 : _issue2_idx_T_59; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_61 = _issue2_idx_T[2] ? 5'h2 : _issue2_idx_T_60; // @[Mux.scala 47:70]
  wire [4:0] _issue2_idx_T_62 = _issue2_idx_T[1] ? 5'h1 : _issue2_idx_T_61; // @[Mux.scala 47:70]
  wire [4:0] issue2_idx = _issue2_idx_T[0] ? 5'h0 : _issue2_idx_T_62; // @[Mux.scala 47:70]
  wire  _issue_num_T = issue1_idx == 5'h1f; // @[reservation_station.scala 87:21]
  wire  _issue_num_T_1 = issue2_idx == 5'h1f; // @[reservation_station.scala 87:53]
  wire  _issue_num_T_2 = issue1_idx == 5'h1f & issue2_idx == 5'h1f; // @[reservation_station.scala 87:40]
  wire  _issue_num_T_4 = issue2_idx != 5'h1f; // @[reservation_station.scala 88:52]
  wire  _issue_num_T_6 = issue1_idx != 5'h1f; // @[reservation_station.scala 88:84]
  wire  _issue_num_T_9 = _issue_num_T & issue2_idx != 5'h1f | issue1_idx != 5'h1f & _issue_num_T_1; // @[reservation_station.scala 88:70]
  wire  _issue_num_T_12 = _issue_num_T_6 & _issue_num_T_4; // @[reservation_station.scala 89:38]
  wire [1:0] _issue_num_T_13 = _issue_num_T_12 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _issue_num_T_14 = _issue_num_T_9 ? 2'h1 : _issue_num_T_13; // @[Mux.scala 101:16]
  wire [1:0] issue_num = _issue_num_T_2 ? 2'h0 : _issue_num_T_14; // @[Mux.scala 101:16]
  wire  _write_num_T = write_idx1 == 5'h1f; // @[reservation_station.scala 98:21]
  wire  _write_num_T_1 = write_idx2 == 5'h1f; // @[reservation_station.scala 98:51]
  wire [31:0] _io_o_issue_packs_0_T_32_pc = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_pc :
    reservation_station_0_io_o_uop_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_32_inst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_inst :
    reservation_station_0_io_o_uop_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_32_func_code = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_func_code :
    reservation_station_0_io_o_uop_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_32_branch_predict_pack_valid = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_valid : reservation_station_0_io_o_uop_branch_predict_pack_valid
    ; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_32_branch_predict_pack_target = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_target :
    reservation_station_0_io_o_uop_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_32_branch_predict_pack_branch_type = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_branch_type :
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_32_branch_predict_pack_select = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_select :
    reservation_station_0_io_o_uop_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_32_branch_predict_pack_taken = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_taken : reservation_station_0_io_o_uop_branch_predict_pack_taken
    ; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_32_phy_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_dst :
    reservation_station_0_io_o_uop_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_32_stale_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_stale_dst :
    reservation_station_0_io_o_uop_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_32_arch_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_dst :
    reservation_station_0_io_o_uop_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_32_inst_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_inst_type :
    reservation_station_0_io_o_uop_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_32_regWen = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_regWen :
    reservation_station_0_io_o_uop_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_32_src1_valid = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src1_valid :
    reservation_station_0_io_o_uop_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_32_phy_rs1 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_rs1 :
    reservation_station_0_io_o_uop_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_32_arch_rs1 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_rs1 :
    reservation_station_0_io_o_uop_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_32_src2_valid = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src2_valid :
    reservation_station_0_io_o_uop_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_32_phy_rs2 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_rs2 :
    reservation_station_0_io_o_uop_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_32_arch_rs2 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_rs2 :
    reservation_station_0_io_o_uop_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_32_rob_idx = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_rob_idx :
    reservation_station_0_io_o_uop_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_32_imm = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_imm :
    reservation_station_0_io_o_uop_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_32_src1_value = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src1_value
     : reservation_station_0_io_o_uop_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_32_src2_value = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src2_value
     : reservation_station_0_io_o_uop_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_32_op1_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_op1_sel :
    reservation_station_0_io_o_uop_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_32_op2_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_op2_sel :
    reservation_station_0_io_o_uop_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_32_alu_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_alu_sel :
    reservation_station_0_io_o_uop_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_32_branch_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_branch_type
     : reservation_station_0_io_o_uop_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_32_mem_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_mem_type :
    reservation_station_0_io_o_uop_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_33_pc = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_pc :
    _io_o_issue_packs_0_T_32_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_33_inst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_inst :
    _io_o_issue_packs_0_T_32_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_33_func_code = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_func_code :
    _io_o_issue_packs_0_T_32_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_33_branch_predict_pack_valid = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_32_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_33_branch_predict_pack_target = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_32_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_33_branch_predict_pack_branch_type = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_32_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_33_branch_predict_pack_select = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_32_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_33_branch_predict_pack_taken = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_32_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_33_phy_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_32_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_33_stale_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_32_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_33_arch_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_32_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_33_inst_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_32_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_33_regWen = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_regWen :
    _io_o_issue_packs_0_T_32_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_33_src1_valid = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_32_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_33_phy_rs1 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_32_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_33_arch_rs1 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_32_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_33_src2_valid = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_32_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_33_phy_rs2 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_32_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_33_arch_rs2 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_32_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_33_rob_idx = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_32_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_33_imm = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_imm :
    _io_o_issue_packs_0_T_32_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_33_src1_value = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_32_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_33_src2_value = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_32_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_33_op1_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_32_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_33_op2_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_32_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_33_alu_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_32_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_33_branch_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_32_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_33_mem_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_32_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_34_pc = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_pc :
    _io_o_issue_packs_0_T_33_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_34_inst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_inst :
    _io_o_issue_packs_0_T_33_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_34_func_code = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_func_code :
    _io_o_issue_packs_0_T_33_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_34_branch_predict_pack_valid = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_33_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_34_branch_predict_pack_target = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_33_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_34_branch_predict_pack_branch_type = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_33_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_34_branch_predict_pack_select = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_33_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_34_branch_predict_pack_taken = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_33_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_34_phy_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_33_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_34_stale_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_33_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_34_arch_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_33_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_34_inst_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_33_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_34_regWen = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_regWen :
    _io_o_issue_packs_0_T_33_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_34_src1_valid = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_33_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_34_phy_rs1 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_33_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_34_arch_rs1 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_33_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_34_src2_valid = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_33_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_34_phy_rs2 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_33_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_34_arch_rs2 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_33_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_34_rob_idx = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_33_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_34_imm = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_imm :
    _io_o_issue_packs_0_T_33_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_34_src1_value = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_33_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_34_src2_value = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_33_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_34_op1_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_33_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_34_op2_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_33_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_34_alu_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_33_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_34_branch_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_33_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_34_mem_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_33_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_35_pc = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_pc :
    _io_o_issue_packs_0_T_34_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_35_inst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_inst :
    _io_o_issue_packs_0_T_34_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_35_func_code = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_func_code :
    _io_o_issue_packs_0_T_34_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_35_branch_predict_pack_valid = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_34_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_35_branch_predict_pack_target = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_34_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_35_branch_predict_pack_branch_type = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_34_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_35_branch_predict_pack_select = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_34_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_35_branch_predict_pack_taken = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_34_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_35_phy_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_34_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_35_stale_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_34_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_35_arch_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_34_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_35_inst_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_34_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_35_regWen = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_regWen :
    _io_o_issue_packs_0_T_34_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_35_src1_valid = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_34_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_35_phy_rs1 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_34_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_35_arch_rs1 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_34_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_35_src2_valid = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_34_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_35_phy_rs2 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_34_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_35_arch_rs2 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_34_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_35_rob_idx = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_34_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_35_imm = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_imm :
    _io_o_issue_packs_0_T_34_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_35_src1_value = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_34_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_35_src2_value = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_34_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_35_op1_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_34_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_35_op2_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_34_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_35_alu_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_34_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_35_branch_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_34_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_35_mem_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_34_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_36_pc = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_pc :
    _io_o_issue_packs_0_T_35_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_36_inst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_inst :
    _io_o_issue_packs_0_T_35_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_36_func_code = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_func_code :
    _io_o_issue_packs_0_T_35_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_36_branch_predict_pack_valid = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_35_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_36_branch_predict_pack_target = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_35_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_36_branch_predict_pack_branch_type = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_35_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_36_branch_predict_pack_select = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_35_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_36_branch_predict_pack_taken = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_35_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_36_phy_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_35_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_36_stale_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_35_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_36_arch_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_35_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_36_inst_type = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_35_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_36_regWen = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_regWen :
    _io_o_issue_packs_0_T_35_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_36_src1_valid = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_35_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_36_phy_rs1 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_35_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_36_arch_rs1 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_35_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_36_src2_valid = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_35_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_36_phy_rs2 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_35_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_36_arch_rs2 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_35_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_36_rob_idx = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_35_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_36_imm = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_imm :
    _io_o_issue_packs_0_T_35_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_36_src1_value = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_35_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_36_src2_value = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_35_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_36_op1_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_35_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_36_op2_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_35_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_36_alu_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_35_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_36_branch_type = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_35_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_36_mem_type = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_35_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_37_pc = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_pc :
    _io_o_issue_packs_0_T_36_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_37_inst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_inst :
    _io_o_issue_packs_0_T_36_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_37_func_code = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_func_code :
    _io_o_issue_packs_0_T_36_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_37_branch_predict_pack_valid = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_36_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_37_branch_predict_pack_target = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_36_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_37_branch_predict_pack_branch_type = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_36_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_37_branch_predict_pack_select = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_36_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_37_branch_predict_pack_taken = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_36_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_37_phy_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_36_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_37_stale_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_36_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_37_arch_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_36_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_37_inst_type = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_36_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_37_regWen = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_regWen :
    _io_o_issue_packs_0_T_36_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_37_src1_valid = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_36_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_37_phy_rs1 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_36_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_37_arch_rs1 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_36_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_37_src2_valid = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_36_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_37_phy_rs2 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_36_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_37_arch_rs2 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_36_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_37_rob_idx = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_36_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_37_imm = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_imm :
    _io_o_issue_packs_0_T_36_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_37_src1_value = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_36_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_37_src2_value = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_36_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_37_op1_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_36_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_37_op2_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_36_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_37_alu_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_36_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_37_branch_type = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_36_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_37_mem_type = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_36_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_38_pc = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_pc :
    _io_o_issue_packs_0_T_37_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_38_inst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_inst :
    _io_o_issue_packs_0_T_37_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_38_func_code = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_func_code :
    _io_o_issue_packs_0_T_37_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_38_branch_predict_pack_valid = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_37_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_38_branch_predict_pack_target = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_37_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_38_branch_predict_pack_branch_type = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_37_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_38_branch_predict_pack_select = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_37_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_38_branch_predict_pack_taken = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_37_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_38_phy_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_37_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_38_stale_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_37_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_38_arch_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_37_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_38_inst_type = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_37_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_38_regWen = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_regWen :
    _io_o_issue_packs_0_T_37_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_38_src1_valid = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_37_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_38_phy_rs1 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_37_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_38_arch_rs1 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_37_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_38_src2_valid = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_37_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_38_phy_rs2 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_37_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_38_arch_rs2 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_37_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_38_rob_idx = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_37_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_38_imm = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_imm :
    _io_o_issue_packs_0_T_37_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_38_src1_value = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_37_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_38_src2_value = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_37_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_38_op1_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_37_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_38_op2_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_37_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_38_alu_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_37_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_38_branch_type = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_37_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_38_mem_type = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_37_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_39_pc = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_pc :
    _io_o_issue_packs_0_T_38_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_39_inst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_inst :
    _io_o_issue_packs_0_T_38_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_39_func_code = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_func_code :
    _io_o_issue_packs_0_T_38_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_39_branch_predict_pack_valid = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_38_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_39_branch_predict_pack_target = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_38_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_39_branch_predict_pack_branch_type = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_38_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_39_branch_predict_pack_select = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_38_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_39_branch_predict_pack_taken = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_38_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_39_phy_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_38_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_39_stale_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_38_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_39_arch_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_38_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_39_inst_type = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_38_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_39_regWen = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_regWen :
    _io_o_issue_packs_0_T_38_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_39_src1_valid = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_38_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_39_phy_rs1 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_38_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_39_arch_rs1 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_38_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_39_src2_valid = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_38_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_39_phy_rs2 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_38_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_39_arch_rs2 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_38_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_39_rob_idx = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_38_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_39_imm = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_imm :
    _io_o_issue_packs_0_T_38_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_39_src1_value = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_38_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_39_src2_value = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_38_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_39_op1_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_38_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_39_op2_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_38_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_39_alu_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_38_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_39_branch_type = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_38_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_39_mem_type = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_38_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_40_pc = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_pc :
    _io_o_issue_packs_0_T_39_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_40_inst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_inst :
    _io_o_issue_packs_0_T_39_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_40_func_code = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_func_code :
    _io_o_issue_packs_0_T_39_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_40_branch_predict_pack_valid = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_39_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_40_branch_predict_pack_target = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_39_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_40_branch_predict_pack_branch_type = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_39_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_40_branch_predict_pack_select = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_39_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_40_branch_predict_pack_taken = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_39_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_40_phy_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_39_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_40_stale_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_39_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_40_arch_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_39_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_40_inst_type = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_39_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_40_regWen = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_regWen :
    _io_o_issue_packs_0_T_39_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_40_src1_valid = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_39_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_40_phy_rs1 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_39_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_40_arch_rs1 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_39_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_40_src2_valid = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_39_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_40_phy_rs2 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_39_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_40_arch_rs2 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_39_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_40_rob_idx = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_39_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_40_imm = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_imm :
    _io_o_issue_packs_0_T_39_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_40_src1_value = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_39_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_40_src2_value = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_39_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_40_op1_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_39_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_40_op2_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_39_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_40_alu_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_39_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_40_branch_type = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_39_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_40_mem_type = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_39_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_41_pc = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_pc :
    _io_o_issue_packs_0_T_40_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_41_inst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_inst :
    _io_o_issue_packs_0_T_40_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_41_func_code = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_func_code :
    _io_o_issue_packs_0_T_40_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_41_branch_predict_pack_valid = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_40_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_41_branch_predict_pack_target = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_40_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_41_branch_predict_pack_branch_type = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_40_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_41_branch_predict_pack_select = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_40_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_41_branch_predict_pack_taken = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_40_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_41_phy_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_40_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_41_stale_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_40_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_41_arch_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_40_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_41_inst_type = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_40_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_41_regWen = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_regWen :
    _io_o_issue_packs_0_T_40_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_41_src1_valid = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_40_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_41_phy_rs1 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_40_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_41_arch_rs1 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_40_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_41_src2_valid = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_40_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_41_phy_rs2 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_40_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_41_arch_rs2 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_40_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_41_rob_idx = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_40_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_41_imm = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_imm :
    _io_o_issue_packs_0_T_40_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_41_src1_value = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_40_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_41_src2_value = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_40_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_41_op1_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_40_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_41_op2_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_40_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_41_alu_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_40_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_41_branch_type = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_40_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_41_mem_type = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_40_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_42_pc = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_pc :
    _io_o_issue_packs_0_T_41_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_42_inst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_inst :
    _io_o_issue_packs_0_T_41_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_42_func_code = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_func_code :
    _io_o_issue_packs_0_T_41_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_42_branch_predict_pack_valid = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_41_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_42_branch_predict_pack_target = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_41_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_42_branch_predict_pack_branch_type = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_41_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_42_branch_predict_pack_select = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_41_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_42_branch_predict_pack_taken = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_41_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_42_phy_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_41_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_42_stale_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_41_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_42_arch_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_41_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_42_inst_type = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_41_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_42_regWen = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_regWen :
    _io_o_issue_packs_0_T_41_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_42_src1_valid = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_41_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_42_phy_rs1 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_41_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_42_arch_rs1 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_41_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_42_src2_valid = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_41_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_42_phy_rs2 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_41_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_42_arch_rs2 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_41_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_42_rob_idx = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_41_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_42_imm = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_imm :
    _io_o_issue_packs_0_T_41_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_42_src1_value = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_41_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_42_src2_value = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_41_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_42_op1_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_41_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_42_op2_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_41_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_42_alu_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_41_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_42_branch_type = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_41_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_42_mem_type = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_41_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_43_pc = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_pc :
    _io_o_issue_packs_0_T_42_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_43_inst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_inst :
    _io_o_issue_packs_0_T_42_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_43_func_code = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_func_code :
    _io_o_issue_packs_0_T_42_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_43_branch_predict_pack_valid = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_42_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_43_branch_predict_pack_target = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_42_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_43_branch_predict_pack_branch_type = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_42_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_43_branch_predict_pack_select = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_42_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_43_branch_predict_pack_taken = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_42_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_43_phy_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_42_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_43_stale_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_42_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_43_arch_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_42_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_43_inst_type = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_42_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_43_regWen = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_regWen :
    _io_o_issue_packs_0_T_42_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_43_src1_valid = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_42_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_43_phy_rs1 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_42_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_43_arch_rs1 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_42_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_43_src2_valid = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_42_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_43_phy_rs2 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_42_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_43_arch_rs2 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_42_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_43_rob_idx = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_42_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_43_imm = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_imm :
    _io_o_issue_packs_0_T_42_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_43_src1_value = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_42_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_43_src2_value = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_42_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_43_op1_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_42_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_43_op2_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_42_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_43_alu_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_42_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_43_branch_type = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_42_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_43_mem_type = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_42_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_44_pc = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_pc :
    _io_o_issue_packs_0_T_43_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_44_inst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_inst :
    _io_o_issue_packs_0_T_43_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_44_func_code = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_func_code :
    _io_o_issue_packs_0_T_43_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_44_branch_predict_pack_valid = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_43_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_44_branch_predict_pack_target = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_43_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_44_branch_predict_pack_branch_type = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_43_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_44_branch_predict_pack_select = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_43_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_44_branch_predict_pack_taken = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_43_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_44_phy_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_43_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_44_stale_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_43_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_44_arch_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_43_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_44_inst_type = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_43_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_44_regWen = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_regWen :
    _io_o_issue_packs_0_T_43_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_44_src1_valid = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_43_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_44_phy_rs1 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_43_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_44_arch_rs1 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_43_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_44_src2_valid = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_43_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_44_phy_rs2 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_43_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_44_arch_rs2 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_43_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_44_rob_idx = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_43_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_44_imm = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_imm :
    _io_o_issue_packs_0_T_43_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_44_src1_value = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_43_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_44_src2_value = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_43_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_44_op1_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_43_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_44_op2_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_43_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_44_alu_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_43_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_44_branch_type = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_43_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_44_mem_type = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_43_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_45_pc = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_pc :
    _io_o_issue_packs_0_T_44_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_45_inst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_inst :
    _io_o_issue_packs_0_T_44_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_45_func_code = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_func_code :
    _io_o_issue_packs_0_T_44_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_45_branch_predict_pack_valid = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_44_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_45_branch_predict_pack_target = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_44_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_45_branch_predict_pack_branch_type = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_44_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_45_branch_predict_pack_select = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_44_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_45_branch_predict_pack_taken = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_44_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_45_phy_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_44_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_45_stale_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_44_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_45_arch_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_44_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_45_inst_type = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_44_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_45_regWen = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_regWen :
    _io_o_issue_packs_0_T_44_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_45_src1_valid = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_44_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_45_phy_rs1 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_44_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_45_arch_rs1 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_44_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_45_src2_valid = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_44_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_45_phy_rs2 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_44_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_45_arch_rs2 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_44_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_45_rob_idx = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_44_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_45_imm = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_imm :
    _io_o_issue_packs_0_T_44_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_45_src1_value = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_44_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_45_src2_value = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_44_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_45_op1_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_44_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_45_op2_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_44_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_45_alu_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_44_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_45_branch_type = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_44_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_45_mem_type = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_44_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_46_pc = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_pc :
    _io_o_issue_packs_0_T_45_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_46_inst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_inst :
    _io_o_issue_packs_0_T_45_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_46_func_code = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_func_code :
    _io_o_issue_packs_0_T_45_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_46_branch_predict_pack_valid = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_45_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_46_branch_predict_pack_target = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_45_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_46_branch_predict_pack_branch_type = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_45_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_46_branch_predict_pack_select = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_45_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_46_branch_predict_pack_taken = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_45_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_46_phy_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_45_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_46_stale_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_45_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_46_arch_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_45_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_46_inst_type = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_45_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_46_regWen = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_regWen :
    _io_o_issue_packs_0_T_45_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_46_src1_valid = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_45_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_46_phy_rs1 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_45_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_46_arch_rs1 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_45_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_46_src2_valid = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_45_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_46_phy_rs2 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_45_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_46_arch_rs2 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_45_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_46_rob_idx = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_45_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_46_imm = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_imm :
    _io_o_issue_packs_0_T_45_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_46_src1_value = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_45_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_46_src2_value = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_45_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_46_op1_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_45_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_46_op2_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_45_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_46_alu_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_45_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_46_branch_type = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_45_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_46_mem_type = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_45_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_47_pc = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_pc :
    _io_o_issue_packs_0_T_46_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_47_inst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_inst :
    _io_o_issue_packs_0_T_46_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_47_func_code = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_func_code :
    _io_o_issue_packs_0_T_46_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_47_branch_predict_pack_valid = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_46_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_47_branch_predict_pack_target = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_46_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_47_branch_predict_pack_branch_type = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_46_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_47_branch_predict_pack_select = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_46_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_47_branch_predict_pack_taken = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_46_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_47_phy_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_46_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_47_stale_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_46_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_47_arch_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_46_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_47_inst_type = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_46_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_47_regWen = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_regWen :
    _io_o_issue_packs_0_T_46_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_47_src1_valid = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_46_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_47_phy_rs1 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_46_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_47_arch_rs1 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_46_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_47_src2_valid = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_46_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_47_phy_rs2 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_46_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_47_arch_rs2 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_46_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_47_rob_idx = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_46_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_47_imm = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_imm :
    _io_o_issue_packs_0_T_46_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_47_src1_value = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_46_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_47_src2_value = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_46_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_47_op1_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_46_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_47_op2_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_46_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_47_alu_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_46_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_47_branch_type = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_46_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_47_mem_type = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_46_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_48_pc = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_pc :
    _io_o_issue_packs_0_T_47_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_48_inst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_inst :
    _io_o_issue_packs_0_T_47_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_48_func_code = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_func_code :
    _io_o_issue_packs_0_T_47_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_48_branch_predict_pack_valid = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_47_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_48_branch_predict_pack_target = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_47_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_48_branch_predict_pack_branch_type = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_47_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_48_branch_predict_pack_select = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_47_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_48_branch_predict_pack_taken = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_47_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_48_phy_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_47_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_48_stale_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_47_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_48_arch_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_47_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_48_inst_type = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_47_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_48_regWen = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_regWen :
    _io_o_issue_packs_0_T_47_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_48_src1_valid = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_47_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_48_phy_rs1 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_47_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_48_arch_rs1 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_47_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_48_src2_valid = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_47_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_48_phy_rs2 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_47_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_48_arch_rs2 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_47_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_48_rob_idx = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_47_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_48_imm = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_imm :
    _io_o_issue_packs_0_T_47_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_48_src1_value = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_47_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_48_src2_value = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_47_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_48_op1_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_47_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_48_op2_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_47_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_48_alu_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_47_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_48_branch_type = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_47_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_48_mem_type = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_47_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_49_pc = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_pc :
    _io_o_issue_packs_0_T_48_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_49_inst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_inst :
    _io_o_issue_packs_0_T_48_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_49_func_code = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_func_code :
    _io_o_issue_packs_0_T_48_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_49_branch_predict_pack_valid = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_48_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_49_branch_predict_pack_target = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_48_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_49_branch_predict_pack_branch_type = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_48_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_49_branch_predict_pack_select = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_48_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_49_branch_predict_pack_taken = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_48_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_49_phy_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_48_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_49_stale_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_48_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_49_arch_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_48_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_49_inst_type = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_48_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_49_regWen = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_regWen :
    _io_o_issue_packs_0_T_48_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_49_src1_valid = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_48_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_49_phy_rs1 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_48_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_49_arch_rs1 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_48_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_49_src2_valid = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_48_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_49_phy_rs2 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_48_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_49_arch_rs2 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_48_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_49_rob_idx = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_48_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_49_imm = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_imm :
    _io_o_issue_packs_0_T_48_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_49_src1_value = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_48_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_49_src2_value = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_48_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_49_op1_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_48_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_49_op2_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_48_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_49_alu_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_48_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_49_branch_type = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_48_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_49_mem_type = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_48_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_50_pc = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_pc :
    _io_o_issue_packs_0_T_49_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_50_inst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_inst :
    _io_o_issue_packs_0_T_49_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_50_func_code = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_func_code :
    _io_o_issue_packs_0_T_49_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_50_branch_predict_pack_valid = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_49_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_50_branch_predict_pack_target = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_49_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_50_branch_predict_pack_branch_type = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_49_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_50_branch_predict_pack_select = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_49_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_50_branch_predict_pack_taken = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_49_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_50_phy_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_49_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_50_stale_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_49_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_50_arch_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_49_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_50_inst_type = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_49_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_50_regWen = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_regWen :
    _io_o_issue_packs_0_T_49_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_50_src1_valid = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_49_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_50_phy_rs1 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_49_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_50_arch_rs1 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_49_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_50_src2_valid = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_49_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_50_phy_rs2 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_49_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_50_arch_rs2 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_49_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_50_rob_idx = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_49_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_50_imm = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_imm :
    _io_o_issue_packs_0_T_49_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_50_src1_value = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_49_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_50_src2_value = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_49_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_50_op1_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_49_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_50_op2_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_49_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_50_alu_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_49_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_50_branch_type = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_49_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_50_mem_type = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_49_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_51_pc = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_pc :
    _io_o_issue_packs_0_T_50_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_51_inst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_inst :
    _io_o_issue_packs_0_T_50_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_51_func_code = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_func_code :
    _io_o_issue_packs_0_T_50_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_51_branch_predict_pack_valid = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_50_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_51_branch_predict_pack_target = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_50_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_51_branch_predict_pack_branch_type = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_50_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_51_branch_predict_pack_select = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_50_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_51_branch_predict_pack_taken = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_50_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_51_phy_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_50_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_51_stale_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_50_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_51_arch_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_50_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_51_inst_type = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_50_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_51_regWen = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_regWen :
    _io_o_issue_packs_0_T_50_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_51_src1_valid = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_50_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_51_phy_rs1 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_50_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_51_arch_rs1 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_50_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_51_src2_valid = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_50_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_51_phy_rs2 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_50_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_51_arch_rs2 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_50_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_51_rob_idx = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_50_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_51_imm = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_imm :
    _io_o_issue_packs_0_T_50_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_51_src1_value = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_50_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_51_src2_value = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_50_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_51_op1_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_50_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_51_op2_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_50_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_51_alu_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_50_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_51_branch_type = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_50_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_51_mem_type = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_50_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_52_pc = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_pc :
    _io_o_issue_packs_0_T_51_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_52_inst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_inst :
    _io_o_issue_packs_0_T_51_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_52_func_code = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_func_code :
    _io_o_issue_packs_0_T_51_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_52_branch_predict_pack_valid = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_51_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_52_branch_predict_pack_target = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_51_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_52_branch_predict_pack_branch_type = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_51_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_52_branch_predict_pack_select = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_51_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_52_branch_predict_pack_taken = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_51_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_52_phy_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_51_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_52_stale_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_51_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_52_arch_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_51_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_52_inst_type = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_51_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_52_regWen = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_regWen :
    _io_o_issue_packs_0_T_51_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_52_src1_valid = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_51_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_52_phy_rs1 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_51_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_52_arch_rs1 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_51_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_52_src2_valid = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_51_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_52_phy_rs2 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_51_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_52_arch_rs2 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_51_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_52_rob_idx = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_51_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_52_imm = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_imm :
    _io_o_issue_packs_0_T_51_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_52_src1_value = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_51_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_52_src2_value = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_51_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_52_op1_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_51_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_52_op2_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_51_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_52_alu_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_51_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_52_branch_type = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_51_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_52_mem_type = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_51_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_53_pc = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_pc :
    _io_o_issue_packs_0_T_52_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_53_inst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_inst :
    _io_o_issue_packs_0_T_52_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_53_func_code = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_func_code :
    _io_o_issue_packs_0_T_52_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_53_branch_predict_pack_valid = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_52_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_53_branch_predict_pack_target = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_52_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_53_branch_predict_pack_branch_type = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_52_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_53_branch_predict_pack_select = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_52_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_53_branch_predict_pack_taken = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_52_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_53_phy_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_52_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_53_stale_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_52_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_53_arch_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_52_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_53_inst_type = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_52_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_53_regWen = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_regWen :
    _io_o_issue_packs_0_T_52_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_53_src1_valid = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_52_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_53_phy_rs1 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_52_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_53_arch_rs1 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_52_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_53_src2_valid = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_52_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_53_phy_rs2 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_52_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_53_arch_rs2 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_52_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_53_rob_idx = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_52_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_53_imm = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_imm :
    _io_o_issue_packs_0_T_52_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_53_src1_value = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_52_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_53_src2_value = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_52_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_53_op1_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_52_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_53_op2_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_52_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_53_alu_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_52_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_53_branch_type = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_52_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_53_mem_type = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_52_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_54_pc = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_pc :
    _io_o_issue_packs_0_T_53_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_54_inst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_inst :
    _io_o_issue_packs_0_T_53_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_54_func_code = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_func_code :
    _io_o_issue_packs_0_T_53_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_54_branch_predict_pack_valid = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_53_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_54_branch_predict_pack_target = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_53_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_54_branch_predict_pack_branch_type = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_53_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_54_branch_predict_pack_select = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_53_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_54_branch_predict_pack_taken = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_53_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_54_phy_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_53_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_54_stale_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_53_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_54_arch_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_53_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_54_inst_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_53_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_54_regWen = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_regWen :
    _io_o_issue_packs_0_T_53_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_54_src1_valid = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_53_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_54_phy_rs1 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_53_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_54_arch_rs1 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_53_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_54_src2_valid = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_53_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_54_phy_rs2 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_53_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_54_arch_rs2 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_53_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_54_rob_idx = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_53_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_54_imm = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_imm :
    _io_o_issue_packs_0_T_53_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_54_src1_value = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_53_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_54_src2_value = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_53_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_54_op1_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_53_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_54_op2_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_53_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_54_alu_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_53_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_54_branch_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_53_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_54_mem_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_53_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_55_pc = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_pc :
    _io_o_issue_packs_0_T_54_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_55_inst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_inst :
    _io_o_issue_packs_0_T_54_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_55_func_code = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_func_code :
    _io_o_issue_packs_0_T_54_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_55_branch_predict_pack_valid = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_54_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_55_branch_predict_pack_target = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_54_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_55_branch_predict_pack_branch_type = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_54_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_55_branch_predict_pack_select = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_54_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_55_branch_predict_pack_taken = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_54_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_55_phy_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_54_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_55_stale_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_54_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_55_arch_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_54_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_55_inst_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_54_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_55_regWen = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_regWen :
    _io_o_issue_packs_0_T_54_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_55_src1_valid = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_54_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_55_phy_rs1 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_54_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_55_arch_rs1 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_54_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_55_src2_valid = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_54_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_55_phy_rs2 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_54_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_55_arch_rs2 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_54_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_55_rob_idx = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_54_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_55_imm = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_imm :
    _io_o_issue_packs_0_T_54_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_55_src1_value = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_54_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_55_src2_value = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_54_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_55_op1_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_54_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_55_op2_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_54_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_55_alu_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_54_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_55_branch_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_54_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_55_mem_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_54_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_56_pc = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_pc :
    _io_o_issue_packs_0_T_55_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_56_inst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_inst :
    _io_o_issue_packs_0_T_55_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_56_func_code = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_func_code :
    _io_o_issue_packs_0_T_55_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_56_branch_predict_pack_valid = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_55_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_56_branch_predict_pack_target = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_55_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_56_branch_predict_pack_branch_type = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_55_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_56_branch_predict_pack_select = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_55_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_56_branch_predict_pack_taken = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_55_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_56_phy_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_55_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_56_stale_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_55_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_56_arch_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_55_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_56_inst_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_55_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_56_regWen = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_regWen :
    _io_o_issue_packs_0_T_55_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_56_src1_valid = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_55_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_56_phy_rs1 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_55_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_56_arch_rs1 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_55_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_56_src2_valid = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_55_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_56_phy_rs2 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_55_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_56_arch_rs2 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_55_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_56_rob_idx = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_55_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_56_imm = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_imm :
    _io_o_issue_packs_0_T_55_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_56_src1_value = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_55_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_56_src2_value = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_55_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_56_op1_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_55_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_56_op2_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_55_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_56_alu_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_55_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_56_branch_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_55_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_56_mem_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_55_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_57_pc = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_pc :
    _io_o_issue_packs_0_T_56_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_57_inst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_inst :
    _io_o_issue_packs_0_T_56_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_57_func_code = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_func_code :
    _io_o_issue_packs_0_T_56_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_57_branch_predict_pack_valid = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_56_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_57_branch_predict_pack_target = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_56_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_57_branch_predict_pack_branch_type = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_56_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_57_branch_predict_pack_select = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_56_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_57_branch_predict_pack_taken = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_56_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_57_phy_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_56_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_57_stale_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_56_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_57_arch_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_56_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_57_inst_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_56_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_57_regWen = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_regWen :
    _io_o_issue_packs_0_T_56_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_57_src1_valid = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_56_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_57_phy_rs1 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_56_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_57_arch_rs1 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_56_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_57_src2_valid = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_56_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_57_phy_rs2 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_56_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_57_arch_rs2 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_56_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_57_rob_idx = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_56_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_57_imm = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_imm :
    _io_o_issue_packs_0_T_56_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_57_src1_value = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_56_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_57_src2_value = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_56_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_57_op1_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_56_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_57_op2_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_56_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_57_alu_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_56_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_57_branch_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_56_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_57_mem_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_56_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_58_pc = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_pc :
    _io_o_issue_packs_0_T_57_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_58_inst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_inst :
    _io_o_issue_packs_0_T_57_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_58_func_code = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_func_code :
    _io_o_issue_packs_0_T_57_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_58_branch_predict_pack_valid = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_57_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_58_branch_predict_pack_target = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_57_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_58_branch_predict_pack_branch_type = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_57_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_58_branch_predict_pack_select = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_57_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_58_branch_predict_pack_taken = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_57_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_58_phy_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_57_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_58_stale_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_57_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_58_arch_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_57_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_58_inst_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_57_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_58_regWen = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_regWen :
    _io_o_issue_packs_0_T_57_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_58_src1_valid = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_57_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_58_phy_rs1 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_57_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_58_arch_rs1 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_57_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_58_src2_valid = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_57_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_58_phy_rs2 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_57_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_58_arch_rs2 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_57_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_58_rob_idx = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_57_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_58_imm = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_imm :
    _io_o_issue_packs_0_T_57_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_58_src1_value = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_57_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_58_src2_value = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_57_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_58_op1_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_57_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_58_op2_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_57_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_58_alu_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_57_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_58_branch_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_57_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_58_mem_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_57_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_59_pc = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_pc :
    _io_o_issue_packs_0_T_58_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_59_inst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_inst :
    _io_o_issue_packs_0_T_58_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_59_func_code = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_func_code :
    _io_o_issue_packs_0_T_58_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_59_branch_predict_pack_valid = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_58_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_59_branch_predict_pack_target = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_58_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_59_branch_predict_pack_branch_type = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_58_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_59_branch_predict_pack_select = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_58_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_59_branch_predict_pack_taken = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_58_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_59_phy_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_58_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_59_stale_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_58_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_59_arch_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_58_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_59_inst_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_58_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_59_regWen = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_regWen :
    _io_o_issue_packs_0_T_58_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_59_src1_valid = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_58_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_59_phy_rs1 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_58_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_59_arch_rs1 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_58_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_59_src2_valid = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_58_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_59_phy_rs2 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_58_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_59_arch_rs2 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_58_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_59_rob_idx = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_58_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_59_imm = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_imm :
    _io_o_issue_packs_0_T_58_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_59_src1_value = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_58_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_59_src2_value = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_58_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_59_op1_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_58_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_59_op2_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_58_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_59_alu_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_58_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_59_branch_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_58_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_59_mem_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_58_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_60_pc = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_pc :
    _io_o_issue_packs_0_T_59_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_60_inst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_inst :
    _io_o_issue_packs_0_T_59_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_60_func_code = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_func_code :
    _io_o_issue_packs_0_T_59_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_60_branch_predict_pack_valid = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_59_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_60_branch_predict_pack_target = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_59_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_60_branch_predict_pack_branch_type = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_59_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_60_branch_predict_pack_select = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_59_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_60_branch_predict_pack_taken = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_59_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_60_phy_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_59_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_60_stale_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_59_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_60_arch_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_59_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_60_inst_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_59_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_60_regWen = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_regWen :
    _io_o_issue_packs_0_T_59_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_60_src1_valid = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_59_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_60_phy_rs1 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_59_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_60_arch_rs1 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_59_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_60_src2_valid = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_59_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_60_phy_rs2 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_59_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_60_arch_rs2 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_59_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_60_rob_idx = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_59_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_60_imm = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_imm :
    _io_o_issue_packs_0_T_59_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_60_src1_value = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_59_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_60_src2_value = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_59_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_60_op1_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_59_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_60_op2_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_59_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_60_alu_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_59_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_60_branch_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_59_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_60_mem_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_59_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_61_pc = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_pc :
    _io_o_issue_packs_0_T_60_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_61_inst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_inst :
    _io_o_issue_packs_0_T_60_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_61_func_code = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_func_code :
    _io_o_issue_packs_0_T_60_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_61_branch_predict_pack_valid = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_60_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_61_branch_predict_pack_target = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_60_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_61_branch_predict_pack_branch_type = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_60_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_61_branch_predict_pack_select = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_60_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_61_branch_predict_pack_taken = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_60_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_61_phy_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_60_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_61_stale_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_60_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_61_arch_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_60_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_61_inst_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_60_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_61_regWen = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_regWen :
    _io_o_issue_packs_0_T_60_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_61_src1_valid = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_60_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_61_phy_rs1 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_60_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_61_arch_rs1 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_60_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_61_src2_valid = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_60_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_61_phy_rs2 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_60_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_61_arch_rs2 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_60_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_61_rob_idx = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_60_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_61_imm = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_imm :
    _io_o_issue_packs_0_T_60_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_61_src1_value = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_60_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_61_src2_value = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_60_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_61_op1_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_60_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_61_op2_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_60_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_61_alu_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_60_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_61_branch_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_60_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_61_mem_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_60_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_62_pc = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_pc :
    _io_o_issue_packs_0_T_61_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_62_inst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_inst :
    _io_o_issue_packs_0_T_61_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_62_func_code = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_func_code :
    _io_o_issue_packs_0_T_61_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_62_branch_predict_pack_valid = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_61_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_62_branch_predict_pack_target = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_61_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_62_branch_predict_pack_branch_type = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_61_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_62_branch_predict_pack_select = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_61_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_62_branch_predict_pack_taken = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_61_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_62_phy_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_61_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_62_stale_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_61_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_62_arch_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_61_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_62_inst_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_61_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_62_regWen = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_regWen :
    _io_o_issue_packs_0_T_61_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_62_src1_valid = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_61_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_62_phy_rs1 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_61_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_62_arch_rs1 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_61_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_62_src2_valid = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_61_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_62_phy_rs2 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_61_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_62_arch_rs2 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_61_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_62_rob_idx = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_61_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_62_imm = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_imm :
    _io_o_issue_packs_0_T_61_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_62_src1_value = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_61_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_62_src2_value = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_61_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_62_op1_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_61_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_62_op2_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_61_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_62_alu_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_61_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_62_branch_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_61_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_62_mem_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_61_mem_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T = 5'h0 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_1 = 5'h1 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_2 = 5'h2 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_3 = 5'h3 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_4 = 5'h4 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_5 = 5'h5 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_6 = 5'h6 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_7 = 5'h7 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_8 = 5'h8 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_9 = 5'h9 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_10 = 5'ha == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_11 = 5'hb == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_12 = 5'hc == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_13 = 5'hd == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_14 = 5'he == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_15 = 5'hf == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_16 = 5'h10 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_17 = 5'h11 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_18 = 5'h12 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_19 = 5'h13 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_20 = 5'h14 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_21 = 5'h15 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_22 = 5'h16 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_23 = 5'h17 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_24 = 5'h18 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_25 = 5'h19 == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_26 = 5'h1a == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_27 = 5'h1b == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_28 = 5'h1c == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_29 = 5'h1d == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_30 = 5'h1e == issue2_idx; // @[reservation_station.scala 107:103]
  wire  _io_o_issue_packs_1_T_31 = 5'h1f == issue2_idx; // @[reservation_station.scala 107:103]
  wire [31:0] _io_o_issue_packs_1_T_32_pc = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_pc :
    reservation_station_0_io_o_uop_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_32_inst = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_inst :
    reservation_station_0_io_o_uop_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_32_func_code = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_func_code
     : reservation_station_0_io_o_uop_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_32_branch_predict_pack_valid = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_valid : reservation_station_0_io_o_uop_branch_predict_pack_valid
    ; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_32_branch_predict_pack_target = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_target :
    reservation_station_0_io_o_uop_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_32_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_branch_type :
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_32_branch_predict_pack_select = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_select :
    reservation_station_0_io_o_uop_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_32_branch_predict_pack_taken = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_taken : reservation_station_0_io_o_uop_branch_predict_pack_taken
    ; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_32_phy_dst = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_phy_dst :
    reservation_station_0_io_o_uop_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_32_stale_dst = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_stale_dst
     : reservation_station_0_io_o_uop_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_32_arch_dst = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_arch_dst :
    reservation_station_0_io_o_uop_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_32_inst_type = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_inst_type
     : reservation_station_0_io_o_uop_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_32_regWen = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_regWen :
    reservation_station_0_io_o_uop_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_32_src1_valid = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_src1_valid :
    reservation_station_0_io_o_uop_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_32_phy_rs1 = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_phy_rs1 :
    reservation_station_0_io_o_uop_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_32_arch_rs1 = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_arch_rs1 :
    reservation_station_0_io_o_uop_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_32_src2_valid = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_src2_valid :
    reservation_station_0_io_o_uop_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_32_phy_rs2 = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_phy_rs2 :
    reservation_station_0_io_o_uop_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_32_arch_rs2 = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_arch_rs2 :
    reservation_station_0_io_o_uop_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_32_rob_idx = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_rob_idx :
    reservation_station_0_io_o_uop_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_32_imm = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_imm :
    reservation_station_0_io_o_uop_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_32_src1_value = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_src1_value : reservation_station_0_io_o_uop_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_32_src2_value = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_src2_value : reservation_station_0_io_o_uop_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_32_op1_sel = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_op1_sel :
    reservation_station_0_io_o_uop_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_32_op2_sel = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_op2_sel :
    reservation_station_0_io_o_uop_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_32_alu_sel = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_alu_sel :
    reservation_station_0_io_o_uop_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_32_branch_type = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_type : reservation_station_0_io_o_uop_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_32_mem_type = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_mem_type :
    reservation_station_0_io_o_uop_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_33_pc = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_pc :
    _io_o_issue_packs_1_T_32_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_33_inst = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_inst :
    _io_o_issue_packs_1_T_32_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_33_func_code = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_func_code
     : _io_o_issue_packs_1_T_32_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_33_branch_predict_pack_valid = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_32_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_33_branch_predict_pack_target = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_32_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_33_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_32_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_33_branch_predict_pack_select = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_32_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_33_branch_predict_pack_taken = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_32_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_33_phy_dst = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_32_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_33_stale_dst = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_32_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_33_arch_dst = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_32_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_33_inst_type = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_32_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_33_regWen = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_regWen :
    _io_o_issue_packs_1_T_32_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_33_src1_valid = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_32_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_33_phy_rs1 = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_32_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_33_arch_rs1 = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_32_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_33_src2_valid = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_32_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_33_phy_rs2 = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_32_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_33_arch_rs2 = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_32_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_33_rob_idx = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_32_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_33_imm = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_imm :
    _io_o_issue_packs_1_T_32_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_33_src1_value = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_src1_value : _io_o_issue_packs_1_T_32_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_33_src2_value = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_src2_value : _io_o_issue_packs_1_T_32_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_33_op1_sel = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_32_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_33_op2_sel = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_32_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_33_alu_sel = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_32_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_33_branch_type = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_type : _io_o_issue_packs_1_T_32_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_33_mem_type = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_32_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_34_pc = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_pc :
    _io_o_issue_packs_1_T_33_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_34_inst = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_inst :
    _io_o_issue_packs_1_T_33_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_34_func_code = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_func_code
     : _io_o_issue_packs_1_T_33_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_34_branch_predict_pack_valid = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_33_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_34_branch_predict_pack_target = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_33_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_34_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_33_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_34_branch_predict_pack_select = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_33_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_34_branch_predict_pack_taken = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_33_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_34_phy_dst = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_33_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_34_stale_dst = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_33_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_34_arch_dst = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_33_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_34_inst_type = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_33_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_34_regWen = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_regWen :
    _io_o_issue_packs_1_T_33_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_34_src1_valid = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_33_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_34_phy_rs1 = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_33_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_34_arch_rs1 = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_33_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_34_src2_valid = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_33_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_34_phy_rs2 = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_33_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_34_arch_rs2 = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_33_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_34_rob_idx = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_33_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_34_imm = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_imm :
    _io_o_issue_packs_1_T_33_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_34_src1_value = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_src1_value : _io_o_issue_packs_1_T_33_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_34_src2_value = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_src2_value : _io_o_issue_packs_1_T_33_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_34_op1_sel = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_33_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_34_op2_sel = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_33_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_34_alu_sel = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_33_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_34_branch_type = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_type : _io_o_issue_packs_1_T_33_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_34_mem_type = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_33_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_35_pc = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_pc :
    _io_o_issue_packs_1_T_34_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_35_inst = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_inst :
    _io_o_issue_packs_1_T_34_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_35_func_code = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_func_code
     : _io_o_issue_packs_1_T_34_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_35_branch_predict_pack_valid = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_34_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_35_branch_predict_pack_target = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_34_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_35_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_34_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_35_branch_predict_pack_select = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_34_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_35_branch_predict_pack_taken = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_34_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_35_phy_dst = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_34_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_35_stale_dst = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_34_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_35_arch_dst = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_34_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_35_inst_type = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_34_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_35_regWen = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_regWen :
    _io_o_issue_packs_1_T_34_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_35_src1_valid = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_34_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_35_phy_rs1 = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_34_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_35_arch_rs1 = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_34_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_35_src2_valid = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_34_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_35_phy_rs2 = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_34_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_35_arch_rs2 = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_34_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_35_rob_idx = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_34_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_35_imm = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_imm :
    _io_o_issue_packs_1_T_34_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_35_src1_value = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_src1_value : _io_o_issue_packs_1_T_34_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_35_src2_value = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_src2_value : _io_o_issue_packs_1_T_34_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_35_op1_sel = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_34_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_35_op2_sel = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_34_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_35_alu_sel = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_34_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_35_branch_type = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_type : _io_o_issue_packs_1_T_34_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_35_mem_type = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_34_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_36_pc = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_pc :
    _io_o_issue_packs_1_T_35_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_36_inst = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_inst :
    _io_o_issue_packs_1_T_35_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_36_func_code = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_func_code
     : _io_o_issue_packs_1_T_35_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_36_branch_predict_pack_valid = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_35_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_36_branch_predict_pack_target = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_35_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_36_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_35_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_36_branch_predict_pack_select = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_35_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_36_branch_predict_pack_taken = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_35_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_36_phy_dst = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_35_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_36_stale_dst = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_35_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_36_arch_dst = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_35_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_36_inst_type = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_35_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_36_regWen = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_regWen :
    _io_o_issue_packs_1_T_35_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_36_src1_valid = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_35_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_36_phy_rs1 = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_35_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_36_arch_rs1 = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_35_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_36_src2_valid = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_35_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_36_phy_rs2 = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_35_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_36_arch_rs2 = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_35_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_36_rob_idx = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_35_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_36_imm = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_imm :
    _io_o_issue_packs_1_T_35_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_36_src1_value = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_src1_value : _io_o_issue_packs_1_T_35_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_36_src2_value = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_src2_value : _io_o_issue_packs_1_T_35_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_36_op1_sel = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_35_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_36_op2_sel = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_35_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_36_alu_sel = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_35_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_36_branch_type = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_type : _io_o_issue_packs_1_T_35_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_36_mem_type = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_35_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_37_pc = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_pc :
    _io_o_issue_packs_1_T_36_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_37_inst = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_inst :
    _io_o_issue_packs_1_T_36_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_37_func_code = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_func_code
     : _io_o_issue_packs_1_T_36_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_37_branch_predict_pack_valid = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_36_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_37_branch_predict_pack_target = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_36_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_37_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_36_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_37_branch_predict_pack_select = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_36_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_37_branch_predict_pack_taken = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_36_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_37_phy_dst = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_36_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_37_stale_dst = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_36_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_37_arch_dst = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_36_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_37_inst_type = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_36_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_37_regWen = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_regWen :
    _io_o_issue_packs_1_T_36_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_37_src1_valid = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_36_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_37_phy_rs1 = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_36_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_37_arch_rs1 = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_36_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_37_src2_valid = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_36_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_37_phy_rs2 = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_36_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_37_arch_rs2 = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_36_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_37_rob_idx = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_36_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_37_imm = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_imm :
    _io_o_issue_packs_1_T_36_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_37_src1_value = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_src1_value : _io_o_issue_packs_1_T_36_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_37_src2_value = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_src2_value : _io_o_issue_packs_1_T_36_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_37_op1_sel = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_36_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_37_op2_sel = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_36_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_37_alu_sel = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_36_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_37_branch_type = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_type : _io_o_issue_packs_1_T_36_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_37_mem_type = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_36_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_38_pc = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_pc :
    _io_o_issue_packs_1_T_37_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_38_inst = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_inst :
    _io_o_issue_packs_1_T_37_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_38_func_code = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_func_code
     : _io_o_issue_packs_1_T_37_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_38_branch_predict_pack_valid = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_37_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_38_branch_predict_pack_target = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_37_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_38_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_37_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_38_branch_predict_pack_select = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_37_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_38_branch_predict_pack_taken = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_37_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_38_phy_dst = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_37_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_38_stale_dst = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_37_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_38_arch_dst = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_37_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_38_inst_type = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_37_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_38_regWen = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_regWen :
    _io_o_issue_packs_1_T_37_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_38_src1_valid = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_37_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_38_phy_rs1 = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_37_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_38_arch_rs1 = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_37_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_38_src2_valid = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_37_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_38_phy_rs2 = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_37_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_38_arch_rs2 = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_37_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_38_rob_idx = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_37_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_38_imm = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_imm :
    _io_o_issue_packs_1_T_37_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_38_src1_value = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_src1_value : _io_o_issue_packs_1_T_37_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_38_src2_value = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_src2_value : _io_o_issue_packs_1_T_37_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_38_op1_sel = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_37_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_38_op2_sel = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_37_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_38_alu_sel = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_37_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_38_branch_type = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_type : _io_o_issue_packs_1_T_37_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_38_mem_type = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_37_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_39_pc = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_pc :
    _io_o_issue_packs_1_T_38_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_39_inst = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_inst :
    _io_o_issue_packs_1_T_38_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_39_func_code = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_func_code
     : _io_o_issue_packs_1_T_38_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_39_branch_predict_pack_valid = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_38_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_39_branch_predict_pack_target = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_38_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_39_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_38_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_39_branch_predict_pack_select = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_38_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_39_branch_predict_pack_taken = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_38_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_39_phy_dst = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_38_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_39_stale_dst = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_38_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_39_arch_dst = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_38_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_39_inst_type = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_38_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_39_regWen = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_regWen :
    _io_o_issue_packs_1_T_38_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_39_src1_valid = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_38_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_39_phy_rs1 = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_38_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_39_arch_rs1 = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_38_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_39_src2_valid = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_38_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_39_phy_rs2 = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_38_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_39_arch_rs2 = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_38_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_39_rob_idx = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_38_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_39_imm = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_imm :
    _io_o_issue_packs_1_T_38_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_39_src1_value = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_src1_value : _io_o_issue_packs_1_T_38_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_39_src2_value = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_src2_value : _io_o_issue_packs_1_T_38_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_39_op1_sel = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_38_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_39_op2_sel = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_38_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_39_alu_sel = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_38_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_39_branch_type = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_type : _io_o_issue_packs_1_T_38_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_39_mem_type = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_38_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_40_pc = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_pc :
    _io_o_issue_packs_1_T_39_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_40_inst = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_inst :
    _io_o_issue_packs_1_T_39_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_40_func_code = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_func_code
     : _io_o_issue_packs_1_T_39_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_40_branch_predict_pack_valid = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_39_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_40_branch_predict_pack_target = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_39_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_40_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_39_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_40_branch_predict_pack_select = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_39_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_40_branch_predict_pack_taken = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_39_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_40_phy_dst = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_39_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_40_stale_dst = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_39_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_40_arch_dst = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_39_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_40_inst_type = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_39_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_40_regWen = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_regWen :
    _io_o_issue_packs_1_T_39_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_40_src1_valid = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_39_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_40_phy_rs1 = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_39_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_40_arch_rs1 = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_39_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_40_src2_valid = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_39_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_40_phy_rs2 = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_39_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_40_arch_rs2 = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_39_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_40_rob_idx = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_39_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_40_imm = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_imm :
    _io_o_issue_packs_1_T_39_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_40_src1_value = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_src1_value : _io_o_issue_packs_1_T_39_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_40_src2_value = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_src2_value : _io_o_issue_packs_1_T_39_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_40_op1_sel = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_39_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_40_op2_sel = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_39_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_40_alu_sel = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_39_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_40_branch_type = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_type : _io_o_issue_packs_1_T_39_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_40_mem_type = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_39_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_41_pc = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_pc :
    _io_o_issue_packs_1_T_40_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_41_inst = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_inst :
    _io_o_issue_packs_1_T_40_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_41_func_code = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_func_code
     : _io_o_issue_packs_1_T_40_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_41_branch_predict_pack_valid = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_40_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_41_branch_predict_pack_target = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_40_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_41_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_40_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_41_branch_predict_pack_select = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_40_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_41_branch_predict_pack_taken = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_40_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_41_phy_dst = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_40_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_41_stale_dst = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_40_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_41_arch_dst = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_40_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_41_inst_type = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_40_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_41_regWen = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_regWen :
    _io_o_issue_packs_1_T_40_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_41_src1_valid = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_40_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_41_phy_rs1 = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_40_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_41_arch_rs1 = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_40_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_41_src2_valid = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_40_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_41_phy_rs2 = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_40_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_41_arch_rs2 = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_40_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_41_rob_idx = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_40_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_41_imm = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_imm :
    _io_o_issue_packs_1_T_40_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_41_src1_value = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_src1_value : _io_o_issue_packs_1_T_40_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_41_src2_value = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_src2_value : _io_o_issue_packs_1_T_40_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_41_op1_sel = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_40_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_41_op2_sel = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_40_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_41_alu_sel = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_40_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_41_branch_type = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_type : _io_o_issue_packs_1_T_40_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_41_mem_type = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_40_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_42_pc = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_pc :
    _io_o_issue_packs_1_T_41_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_42_inst = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_inst :
    _io_o_issue_packs_1_T_41_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_42_func_code = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_func_code
     : _io_o_issue_packs_1_T_41_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_42_branch_predict_pack_valid = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_41_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_42_branch_predict_pack_target = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_41_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_42_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_41_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_42_branch_predict_pack_select = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_41_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_42_branch_predict_pack_taken = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_41_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_42_phy_dst = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_41_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_42_stale_dst = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_41_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_42_arch_dst = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_41_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_42_inst_type = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_41_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_42_regWen = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_regWen :
    _io_o_issue_packs_1_T_41_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_42_src1_valid = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_41_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_42_phy_rs1 = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_41_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_42_arch_rs1 = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_41_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_42_src2_valid = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_41_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_42_phy_rs2 = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_41_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_42_arch_rs2 = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_41_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_42_rob_idx = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_41_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_42_imm = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_imm :
    _io_o_issue_packs_1_T_41_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_42_src1_value = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_src1_value : _io_o_issue_packs_1_T_41_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_42_src2_value = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_src2_value : _io_o_issue_packs_1_T_41_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_42_op1_sel = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_41_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_42_op2_sel = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_41_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_42_alu_sel = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_41_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_42_branch_type = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_type : _io_o_issue_packs_1_T_41_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_42_mem_type = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_41_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_43_pc = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_pc :
    _io_o_issue_packs_1_T_42_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_43_inst = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_inst :
    _io_o_issue_packs_1_T_42_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_43_func_code = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_func_code
     : _io_o_issue_packs_1_T_42_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_43_branch_predict_pack_valid = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_42_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_43_branch_predict_pack_target = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_42_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_43_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_42_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_43_branch_predict_pack_select = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_42_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_43_branch_predict_pack_taken = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_42_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_43_phy_dst = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_42_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_43_stale_dst = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_42_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_43_arch_dst = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_42_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_43_inst_type = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_42_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_43_regWen = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_regWen :
    _io_o_issue_packs_1_T_42_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_43_src1_valid = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_42_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_43_phy_rs1 = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_42_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_43_arch_rs1 = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_42_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_43_src2_valid = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_42_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_43_phy_rs2 = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_42_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_43_arch_rs2 = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_42_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_43_rob_idx = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_42_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_43_imm = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_imm :
    _io_o_issue_packs_1_T_42_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_43_src1_value = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_src1_value : _io_o_issue_packs_1_T_42_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_43_src2_value = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_src2_value : _io_o_issue_packs_1_T_42_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_43_op1_sel = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_42_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_43_op2_sel = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_42_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_43_alu_sel = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_42_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_43_branch_type = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_type : _io_o_issue_packs_1_T_42_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_43_mem_type = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_42_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_44_pc = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_pc :
    _io_o_issue_packs_1_T_43_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_44_inst = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_inst :
    _io_o_issue_packs_1_T_43_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_44_func_code = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_func_code
     : _io_o_issue_packs_1_T_43_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_44_branch_predict_pack_valid = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_43_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_44_branch_predict_pack_target = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_43_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_44_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_43_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_44_branch_predict_pack_select = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_43_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_44_branch_predict_pack_taken = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_43_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_44_phy_dst = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_43_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_44_stale_dst = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_43_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_44_arch_dst = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_43_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_44_inst_type = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_43_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_44_regWen = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_regWen :
    _io_o_issue_packs_1_T_43_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_44_src1_valid = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_43_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_44_phy_rs1 = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_43_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_44_arch_rs1 = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_43_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_44_src2_valid = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_43_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_44_phy_rs2 = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_43_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_44_arch_rs2 = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_43_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_44_rob_idx = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_43_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_44_imm = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_imm :
    _io_o_issue_packs_1_T_43_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_44_src1_value = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_src1_value : _io_o_issue_packs_1_T_43_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_44_src2_value = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_src2_value : _io_o_issue_packs_1_T_43_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_44_op1_sel = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_43_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_44_op2_sel = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_43_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_44_alu_sel = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_43_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_44_branch_type = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_type : _io_o_issue_packs_1_T_43_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_44_mem_type = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_43_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_45_pc = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_pc :
    _io_o_issue_packs_1_T_44_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_45_inst = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_inst :
    _io_o_issue_packs_1_T_44_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_45_func_code = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_func_code
     : _io_o_issue_packs_1_T_44_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_45_branch_predict_pack_valid = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_44_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_45_branch_predict_pack_target = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_44_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_45_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_44_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_45_branch_predict_pack_select = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_44_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_45_branch_predict_pack_taken = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_44_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_45_phy_dst = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_44_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_45_stale_dst = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_44_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_45_arch_dst = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_44_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_45_inst_type = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_44_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_45_regWen = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_regWen :
    _io_o_issue_packs_1_T_44_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_45_src1_valid = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_44_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_45_phy_rs1 = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_44_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_45_arch_rs1 = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_44_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_45_src2_valid = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_44_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_45_phy_rs2 = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_44_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_45_arch_rs2 = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_44_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_45_rob_idx = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_44_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_45_imm = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_imm :
    _io_o_issue_packs_1_T_44_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_45_src1_value = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_src1_value : _io_o_issue_packs_1_T_44_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_45_src2_value = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_src2_value : _io_o_issue_packs_1_T_44_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_45_op1_sel = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_44_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_45_op2_sel = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_44_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_45_alu_sel = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_44_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_45_branch_type = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_type : _io_o_issue_packs_1_T_44_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_45_mem_type = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_44_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_46_pc = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_pc :
    _io_o_issue_packs_1_T_45_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_46_inst = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_inst :
    _io_o_issue_packs_1_T_45_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_46_func_code = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_func_code
     : _io_o_issue_packs_1_T_45_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_46_branch_predict_pack_valid = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_45_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_46_branch_predict_pack_target = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_45_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_46_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_45_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_46_branch_predict_pack_select = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_45_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_46_branch_predict_pack_taken = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_45_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_46_phy_dst = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_45_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_46_stale_dst = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_45_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_46_arch_dst = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_45_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_46_inst_type = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_45_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_46_regWen = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_regWen :
    _io_o_issue_packs_1_T_45_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_46_src1_valid = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_45_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_46_phy_rs1 = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_45_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_46_arch_rs1 = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_45_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_46_src2_valid = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_45_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_46_phy_rs2 = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_45_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_46_arch_rs2 = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_45_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_46_rob_idx = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_45_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_46_imm = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_imm :
    _io_o_issue_packs_1_T_45_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_46_src1_value = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_src1_value : _io_o_issue_packs_1_T_45_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_46_src2_value = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_src2_value : _io_o_issue_packs_1_T_45_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_46_op1_sel = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_45_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_46_op2_sel = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_45_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_46_alu_sel = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_45_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_46_branch_type = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_type : _io_o_issue_packs_1_T_45_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_46_mem_type = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_45_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_47_pc = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_pc :
    _io_o_issue_packs_1_T_46_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_47_inst = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_inst :
    _io_o_issue_packs_1_T_46_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_47_func_code = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_func_code
     : _io_o_issue_packs_1_T_46_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_47_branch_predict_pack_valid = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_46_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_47_branch_predict_pack_target = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_46_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_47_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_46_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_47_branch_predict_pack_select = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_46_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_47_branch_predict_pack_taken = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_46_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_47_phy_dst = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_46_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_47_stale_dst = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_46_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_47_arch_dst = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_46_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_47_inst_type = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_46_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_47_regWen = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_regWen :
    _io_o_issue_packs_1_T_46_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_47_src1_valid = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_46_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_47_phy_rs1 = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_46_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_47_arch_rs1 = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_46_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_47_src2_valid = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_46_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_47_phy_rs2 = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_46_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_47_arch_rs2 = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_46_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_47_rob_idx = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_46_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_47_imm = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_imm :
    _io_o_issue_packs_1_T_46_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_47_src1_value = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_src1_value : _io_o_issue_packs_1_T_46_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_47_src2_value = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_src2_value : _io_o_issue_packs_1_T_46_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_47_op1_sel = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_46_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_47_op2_sel = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_46_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_47_alu_sel = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_46_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_47_branch_type = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_type : _io_o_issue_packs_1_T_46_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_47_mem_type = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_46_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_48_pc = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_pc :
    _io_o_issue_packs_1_T_47_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_48_inst = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_inst :
    _io_o_issue_packs_1_T_47_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_48_func_code = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_func_code
     : _io_o_issue_packs_1_T_47_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_48_branch_predict_pack_valid = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_47_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_48_branch_predict_pack_target = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_47_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_48_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_47_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_48_branch_predict_pack_select = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_47_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_48_branch_predict_pack_taken = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_47_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_48_phy_dst = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_47_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_48_stale_dst = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_47_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_48_arch_dst = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_47_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_48_inst_type = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_47_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_48_regWen = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_regWen :
    _io_o_issue_packs_1_T_47_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_48_src1_valid = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_47_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_48_phy_rs1 = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_47_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_48_arch_rs1 = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_47_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_48_src2_valid = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_47_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_48_phy_rs2 = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_47_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_48_arch_rs2 = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_47_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_48_rob_idx = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_47_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_48_imm = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_imm :
    _io_o_issue_packs_1_T_47_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_48_src1_value = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_src1_value : _io_o_issue_packs_1_T_47_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_48_src2_value = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_src2_value : _io_o_issue_packs_1_T_47_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_48_op1_sel = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_47_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_48_op2_sel = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_47_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_48_alu_sel = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_47_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_48_branch_type = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_type : _io_o_issue_packs_1_T_47_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_48_mem_type = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_47_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_49_pc = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_pc :
    _io_o_issue_packs_1_T_48_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_49_inst = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_inst :
    _io_o_issue_packs_1_T_48_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_49_func_code = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_func_code
     : _io_o_issue_packs_1_T_48_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_49_branch_predict_pack_valid = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_48_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_49_branch_predict_pack_target = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_48_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_49_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_48_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_49_branch_predict_pack_select = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_48_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_49_branch_predict_pack_taken = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_48_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_49_phy_dst = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_48_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_49_stale_dst = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_48_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_49_arch_dst = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_48_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_49_inst_type = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_48_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_49_regWen = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_regWen :
    _io_o_issue_packs_1_T_48_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_49_src1_valid = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_48_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_49_phy_rs1 = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_48_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_49_arch_rs1 = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_48_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_49_src2_valid = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_48_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_49_phy_rs2 = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_48_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_49_arch_rs2 = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_48_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_49_rob_idx = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_48_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_49_imm = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_imm :
    _io_o_issue_packs_1_T_48_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_49_src1_value = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_src1_value : _io_o_issue_packs_1_T_48_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_49_src2_value = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_src2_value : _io_o_issue_packs_1_T_48_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_49_op1_sel = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_48_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_49_op2_sel = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_48_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_49_alu_sel = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_48_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_49_branch_type = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_type : _io_o_issue_packs_1_T_48_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_49_mem_type = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_48_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_50_pc = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_pc :
    _io_o_issue_packs_1_T_49_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_50_inst = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_inst :
    _io_o_issue_packs_1_T_49_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_50_func_code = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_func_code
     : _io_o_issue_packs_1_T_49_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_50_branch_predict_pack_valid = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_49_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_50_branch_predict_pack_target = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_49_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_50_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_49_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_50_branch_predict_pack_select = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_49_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_50_branch_predict_pack_taken = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_49_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_50_phy_dst = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_49_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_50_stale_dst = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_49_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_50_arch_dst = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_49_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_50_inst_type = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_49_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_50_regWen = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_regWen :
    _io_o_issue_packs_1_T_49_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_50_src1_valid = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_49_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_50_phy_rs1 = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_49_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_50_arch_rs1 = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_49_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_50_src2_valid = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_49_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_50_phy_rs2 = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_49_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_50_arch_rs2 = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_49_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_50_rob_idx = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_49_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_50_imm = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_imm :
    _io_o_issue_packs_1_T_49_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_50_src1_value = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_src1_value : _io_o_issue_packs_1_T_49_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_50_src2_value = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_src2_value : _io_o_issue_packs_1_T_49_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_50_op1_sel = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_49_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_50_op2_sel = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_49_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_50_alu_sel = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_49_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_50_branch_type = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_type : _io_o_issue_packs_1_T_49_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_50_mem_type = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_49_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_51_pc = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_pc :
    _io_o_issue_packs_1_T_50_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_51_inst = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_inst :
    _io_o_issue_packs_1_T_50_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_51_func_code = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_func_code
     : _io_o_issue_packs_1_T_50_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_51_branch_predict_pack_valid = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_50_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_51_branch_predict_pack_target = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_50_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_51_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_50_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_51_branch_predict_pack_select = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_50_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_51_branch_predict_pack_taken = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_50_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_51_phy_dst = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_50_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_51_stale_dst = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_50_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_51_arch_dst = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_50_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_51_inst_type = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_50_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_51_regWen = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_regWen :
    _io_o_issue_packs_1_T_50_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_51_src1_valid = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_50_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_51_phy_rs1 = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_50_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_51_arch_rs1 = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_50_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_51_src2_valid = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_50_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_51_phy_rs2 = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_50_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_51_arch_rs2 = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_50_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_51_rob_idx = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_50_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_51_imm = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_imm :
    _io_o_issue_packs_1_T_50_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_51_src1_value = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_src1_value : _io_o_issue_packs_1_T_50_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_51_src2_value = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_src2_value : _io_o_issue_packs_1_T_50_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_51_op1_sel = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_50_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_51_op2_sel = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_50_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_51_alu_sel = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_50_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_51_branch_type = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_type : _io_o_issue_packs_1_T_50_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_51_mem_type = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_50_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_52_pc = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_pc :
    _io_o_issue_packs_1_T_51_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_52_inst = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_inst :
    _io_o_issue_packs_1_T_51_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_52_func_code = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_func_code
     : _io_o_issue_packs_1_T_51_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_52_branch_predict_pack_valid = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_51_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_52_branch_predict_pack_target = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_51_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_52_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_51_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_52_branch_predict_pack_select = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_51_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_52_branch_predict_pack_taken = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_51_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_52_phy_dst = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_51_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_52_stale_dst = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_51_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_52_arch_dst = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_51_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_52_inst_type = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_51_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_52_regWen = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_regWen :
    _io_o_issue_packs_1_T_51_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_52_src1_valid = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_51_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_52_phy_rs1 = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_51_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_52_arch_rs1 = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_51_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_52_src2_valid = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_51_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_52_phy_rs2 = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_51_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_52_arch_rs2 = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_51_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_52_rob_idx = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_51_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_52_imm = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_imm :
    _io_o_issue_packs_1_T_51_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_52_src1_value = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_src1_value : _io_o_issue_packs_1_T_51_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_52_src2_value = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_src2_value : _io_o_issue_packs_1_T_51_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_52_op1_sel = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_51_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_52_op2_sel = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_51_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_52_alu_sel = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_51_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_52_branch_type = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_type : _io_o_issue_packs_1_T_51_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_52_mem_type = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_51_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_53_pc = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_pc :
    _io_o_issue_packs_1_T_52_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_53_inst = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_inst :
    _io_o_issue_packs_1_T_52_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_53_func_code = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_func_code
     : _io_o_issue_packs_1_T_52_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_53_branch_predict_pack_valid = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_52_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_53_branch_predict_pack_target = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_52_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_53_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_52_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_53_branch_predict_pack_select = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_52_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_53_branch_predict_pack_taken = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_52_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_53_phy_dst = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_52_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_53_stale_dst = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_52_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_53_arch_dst = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_52_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_53_inst_type = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_52_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_53_regWen = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_regWen :
    _io_o_issue_packs_1_T_52_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_53_src1_valid = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_52_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_53_phy_rs1 = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_52_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_53_arch_rs1 = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_52_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_53_src2_valid = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_52_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_53_phy_rs2 = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_52_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_53_arch_rs2 = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_52_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_53_rob_idx = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_52_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_53_imm = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_imm :
    _io_o_issue_packs_1_T_52_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_53_src1_value = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_src1_value : _io_o_issue_packs_1_T_52_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_53_src2_value = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_src2_value : _io_o_issue_packs_1_T_52_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_53_op1_sel = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_52_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_53_op2_sel = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_52_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_53_alu_sel = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_52_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_53_branch_type = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_type : _io_o_issue_packs_1_T_52_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_53_mem_type = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_52_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_54_pc = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_pc :
    _io_o_issue_packs_1_T_53_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_54_inst = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_inst :
    _io_o_issue_packs_1_T_53_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_54_func_code = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_func_code :
    _io_o_issue_packs_1_T_53_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_54_branch_predict_pack_valid = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_53_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_54_branch_predict_pack_target = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_53_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_54_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_53_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_54_branch_predict_pack_select = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_53_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_54_branch_predict_pack_taken = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_53_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_54_phy_dst = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_53_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_54_stale_dst = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_53_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_54_arch_dst = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_53_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_54_inst_type = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_53_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_54_regWen = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_regWen :
    _io_o_issue_packs_1_T_53_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_54_src1_valid = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_53_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_54_phy_rs1 = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_53_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_54_arch_rs1 = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_53_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_54_src2_valid = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_53_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_54_phy_rs2 = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_53_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_54_arch_rs2 = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_53_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_54_rob_idx = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_53_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_54_imm = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_imm :
    _io_o_issue_packs_1_T_53_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_54_src1_value = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_53_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_54_src2_value = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_53_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_54_op1_sel = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_53_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_54_op2_sel = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_53_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_54_alu_sel = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_53_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_54_branch_type = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_53_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_54_mem_type = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_53_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_55_pc = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_pc :
    _io_o_issue_packs_1_T_54_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_55_inst = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_inst :
    _io_o_issue_packs_1_T_54_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_55_func_code = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_func_code :
    _io_o_issue_packs_1_T_54_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_55_branch_predict_pack_valid = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_54_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_55_branch_predict_pack_target = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_54_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_55_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_54_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_55_branch_predict_pack_select = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_54_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_55_branch_predict_pack_taken = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_54_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_55_phy_dst = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_54_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_55_stale_dst = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_54_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_55_arch_dst = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_54_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_55_inst_type = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_54_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_55_regWen = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_regWen :
    _io_o_issue_packs_1_T_54_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_55_src1_valid = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_54_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_55_phy_rs1 = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_54_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_55_arch_rs1 = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_54_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_55_src2_valid = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_54_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_55_phy_rs2 = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_54_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_55_arch_rs2 = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_54_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_55_rob_idx = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_54_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_55_imm = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_imm :
    _io_o_issue_packs_1_T_54_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_55_src1_value = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_54_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_55_src2_value = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_54_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_55_op1_sel = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_54_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_55_op2_sel = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_54_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_55_alu_sel = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_54_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_55_branch_type = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_54_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_55_mem_type = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_54_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_56_pc = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_pc :
    _io_o_issue_packs_1_T_55_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_56_inst = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_inst :
    _io_o_issue_packs_1_T_55_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_56_func_code = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_func_code :
    _io_o_issue_packs_1_T_55_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_56_branch_predict_pack_valid = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_55_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_56_branch_predict_pack_target = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_55_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_56_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_55_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_56_branch_predict_pack_select = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_55_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_56_branch_predict_pack_taken = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_55_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_56_phy_dst = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_55_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_56_stale_dst = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_55_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_56_arch_dst = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_55_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_56_inst_type = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_55_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_56_regWen = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_regWen :
    _io_o_issue_packs_1_T_55_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_56_src1_valid = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_55_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_56_phy_rs1 = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_55_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_56_arch_rs1 = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_55_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_56_src2_valid = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_55_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_56_phy_rs2 = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_55_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_56_arch_rs2 = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_55_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_56_rob_idx = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_55_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_56_imm = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_imm :
    _io_o_issue_packs_1_T_55_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_56_src1_value = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_55_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_56_src2_value = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_55_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_56_op1_sel = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_55_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_56_op2_sel = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_55_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_56_alu_sel = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_55_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_56_branch_type = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_55_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_56_mem_type = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_55_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_57_pc = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_pc :
    _io_o_issue_packs_1_T_56_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_57_inst = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_inst :
    _io_o_issue_packs_1_T_56_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_57_func_code = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_func_code :
    _io_o_issue_packs_1_T_56_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_57_branch_predict_pack_valid = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_56_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_57_branch_predict_pack_target = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_56_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_57_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_56_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_57_branch_predict_pack_select = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_56_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_57_branch_predict_pack_taken = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_56_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_57_phy_dst = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_56_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_57_stale_dst = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_56_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_57_arch_dst = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_56_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_57_inst_type = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_56_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_57_regWen = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_regWen :
    _io_o_issue_packs_1_T_56_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_57_src1_valid = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_56_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_57_phy_rs1 = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_56_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_57_arch_rs1 = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_56_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_57_src2_valid = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_56_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_57_phy_rs2 = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_56_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_57_arch_rs2 = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_56_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_57_rob_idx = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_56_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_57_imm = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_imm :
    _io_o_issue_packs_1_T_56_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_57_src1_value = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_56_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_57_src2_value = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_56_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_57_op1_sel = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_56_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_57_op2_sel = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_56_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_57_alu_sel = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_56_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_57_branch_type = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_56_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_57_mem_type = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_56_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_58_pc = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_pc :
    _io_o_issue_packs_1_T_57_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_58_inst = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_inst :
    _io_o_issue_packs_1_T_57_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_58_func_code = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_func_code :
    _io_o_issue_packs_1_T_57_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_58_branch_predict_pack_valid = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_57_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_58_branch_predict_pack_target = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_57_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_58_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_57_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_58_branch_predict_pack_select = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_57_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_58_branch_predict_pack_taken = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_57_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_58_phy_dst = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_57_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_58_stale_dst = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_57_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_58_arch_dst = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_57_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_58_inst_type = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_57_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_58_regWen = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_regWen :
    _io_o_issue_packs_1_T_57_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_58_src1_valid = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_57_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_58_phy_rs1 = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_57_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_58_arch_rs1 = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_57_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_58_src2_valid = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_57_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_58_phy_rs2 = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_57_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_58_arch_rs2 = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_57_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_58_rob_idx = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_57_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_58_imm = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_imm :
    _io_o_issue_packs_1_T_57_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_58_src1_value = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_57_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_58_src2_value = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_57_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_58_op1_sel = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_57_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_58_op2_sel = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_57_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_58_alu_sel = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_57_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_58_branch_type = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_57_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_58_mem_type = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_57_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_59_pc = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_pc :
    _io_o_issue_packs_1_T_58_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_59_inst = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_inst :
    _io_o_issue_packs_1_T_58_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_59_func_code = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_func_code :
    _io_o_issue_packs_1_T_58_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_59_branch_predict_pack_valid = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_58_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_59_branch_predict_pack_target = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_58_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_59_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_58_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_59_branch_predict_pack_select = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_58_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_59_branch_predict_pack_taken = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_58_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_59_phy_dst = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_58_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_59_stale_dst = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_58_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_59_arch_dst = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_58_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_59_inst_type = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_58_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_59_regWen = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_regWen :
    _io_o_issue_packs_1_T_58_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_59_src1_valid = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_58_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_59_phy_rs1 = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_58_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_59_arch_rs1 = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_58_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_59_src2_valid = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_58_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_59_phy_rs2 = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_58_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_59_arch_rs2 = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_58_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_59_rob_idx = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_58_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_59_imm = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_imm :
    _io_o_issue_packs_1_T_58_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_59_src1_value = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_58_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_59_src2_value = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_58_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_59_op1_sel = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_58_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_59_op2_sel = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_58_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_59_alu_sel = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_58_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_59_branch_type = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_58_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_59_mem_type = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_58_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_60_pc = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_pc :
    _io_o_issue_packs_1_T_59_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_60_inst = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_inst :
    _io_o_issue_packs_1_T_59_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_60_func_code = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_func_code :
    _io_o_issue_packs_1_T_59_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_60_branch_predict_pack_valid = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_59_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_60_branch_predict_pack_target = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_59_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_60_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_59_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_60_branch_predict_pack_select = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_59_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_60_branch_predict_pack_taken = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_59_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_60_phy_dst = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_59_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_60_stale_dst = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_59_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_60_arch_dst = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_59_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_60_inst_type = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_59_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_60_regWen = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_regWen :
    _io_o_issue_packs_1_T_59_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_60_src1_valid = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_59_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_60_phy_rs1 = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_59_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_60_arch_rs1 = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_59_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_60_src2_valid = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_59_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_60_phy_rs2 = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_59_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_60_arch_rs2 = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_59_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_60_rob_idx = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_59_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_60_imm = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_imm :
    _io_o_issue_packs_1_T_59_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_60_src1_value = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_59_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_60_src2_value = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_59_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_60_op1_sel = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_59_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_60_op2_sel = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_59_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_60_alu_sel = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_59_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_60_branch_type = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_59_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_60_mem_type = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_59_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_61_pc = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_pc :
    _io_o_issue_packs_1_T_60_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_61_inst = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_inst :
    _io_o_issue_packs_1_T_60_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_61_func_code = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_func_code :
    _io_o_issue_packs_1_T_60_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_61_branch_predict_pack_valid = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_60_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_61_branch_predict_pack_target = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_60_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_61_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_60_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_61_branch_predict_pack_select = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_60_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_61_branch_predict_pack_taken = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_60_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_61_phy_dst = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_60_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_61_stale_dst = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_60_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_61_arch_dst = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_60_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_61_inst_type = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_60_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_61_regWen = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_regWen :
    _io_o_issue_packs_1_T_60_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_61_src1_valid = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_60_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_61_phy_rs1 = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_60_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_61_arch_rs1 = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_60_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_61_src2_valid = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_60_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_61_phy_rs2 = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_60_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_61_arch_rs2 = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_60_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_61_rob_idx = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_60_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_61_imm = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_imm :
    _io_o_issue_packs_1_T_60_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_61_src1_value = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_60_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_61_src2_value = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_60_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_61_op1_sel = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_60_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_61_op2_sel = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_60_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_61_alu_sel = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_60_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_61_branch_type = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_60_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_61_mem_type = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_60_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_62_pc = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_pc :
    _io_o_issue_packs_1_T_61_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_62_inst = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_inst :
    _io_o_issue_packs_1_T_61_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_62_func_code = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_func_code :
    _io_o_issue_packs_1_T_61_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_62_branch_predict_pack_valid = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_61_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_62_branch_predict_pack_target = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_61_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_62_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_61_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_62_branch_predict_pack_select = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_61_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_62_branch_predict_pack_taken = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_61_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_62_phy_dst = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_61_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_62_stale_dst = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_61_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_62_arch_dst = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_61_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_62_inst_type = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_61_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_62_regWen = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_regWen :
    _io_o_issue_packs_1_T_61_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_62_src1_valid = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_61_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_62_phy_rs1 = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_61_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_62_arch_rs1 = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_61_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_62_src2_valid = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_61_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_62_phy_rs2 = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_61_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_62_arch_rs2 = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_61_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_62_rob_idx = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_61_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_62_imm = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_imm :
    _io_o_issue_packs_1_T_61_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_62_src1_value = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_61_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_62_src2_value = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_61_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_62_op1_sel = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_61_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_62_op2_sel = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_61_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_62_alu_sel = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_61_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_62_branch_type = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_61_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_62_mem_type = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_61_mem_type; // @[Mux.scala 101:16]
  wire  _reservation_station_0_io_i_write_slot_T = 5'h0 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_0_io_i_write_slot_T_2 = 5'h0 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_0_io_i_write_slot_T_5 = 5'h0 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_1_io_i_write_slot_T = 5'h1 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_1_io_i_write_slot_T_2 = 5'h1 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_1_io_i_write_slot_T_5 = 5'h1 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_2_io_i_write_slot_T = 5'h2 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_2_io_i_write_slot_T_2 = 5'h2 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_2_io_i_write_slot_T_5 = 5'h2 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_3_io_i_write_slot_T = 5'h3 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_3_io_i_write_slot_T_2 = 5'h3 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_3_io_i_write_slot_T_5 = 5'h3 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_4_io_i_write_slot_T = 5'h4 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_4_io_i_write_slot_T_2 = 5'h4 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_4_io_i_write_slot_T_5 = 5'h4 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_5_io_i_write_slot_T = 5'h5 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_5_io_i_write_slot_T_2 = 5'h5 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_5_io_i_write_slot_T_5 = 5'h5 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_6_io_i_write_slot_T = 5'h6 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_6_io_i_write_slot_T_2 = 5'h6 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_6_io_i_write_slot_T_5 = 5'h6 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_7_io_i_write_slot_T = 5'h7 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_7_io_i_write_slot_T_2 = 5'h7 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_7_io_i_write_slot_T_5 = 5'h7 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_8_io_i_write_slot_T = 5'h8 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_8_io_i_write_slot_T_2 = 5'h8 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_8_io_i_write_slot_T_5 = 5'h8 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_9_io_i_write_slot_T = 5'h9 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_9_io_i_write_slot_T_2 = 5'h9 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_9_io_i_write_slot_T_5 = 5'h9 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_10_io_i_write_slot_T = 5'ha == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_10_io_i_write_slot_T_2 = 5'ha == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_10_io_i_write_slot_T_5 = 5'ha == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_11_io_i_write_slot_T = 5'hb == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_11_io_i_write_slot_T_2 = 5'hb == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_11_io_i_write_slot_T_5 = 5'hb == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_12_io_i_write_slot_T = 5'hc == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_12_io_i_write_slot_T_2 = 5'hc == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_12_io_i_write_slot_T_5 = 5'hc == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_13_io_i_write_slot_T = 5'hd == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_13_io_i_write_slot_T_2 = 5'hd == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_13_io_i_write_slot_T_5 = 5'hd == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_14_io_i_write_slot_T = 5'he == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_14_io_i_write_slot_T_2 = 5'he == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_14_io_i_write_slot_T_5 = 5'he == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_15_io_i_write_slot_T = 5'hf == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_15_io_i_write_slot_T_2 = 5'hf == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_15_io_i_write_slot_T_5 = 5'hf == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_16_io_i_write_slot_T = 5'h10 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_16_io_i_write_slot_T_2 = 5'h10 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_16_io_i_write_slot_T_5 = 5'h10 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_17_io_i_write_slot_T = 5'h11 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_17_io_i_write_slot_T_2 = 5'h11 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_17_io_i_write_slot_T_5 = 5'h11 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_18_io_i_write_slot_T = 5'h12 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_18_io_i_write_slot_T_2 = 5'h12 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_18_io_i_write_slot_T_5 = 5'h12 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_19_io_i_write_slot_T = 5'h13 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_19_io_i_write_slot_T_2 = 5'h13 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_19_io_i_write_slot_T_5 = 5'h13 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_20_io_i_write_slot_T = 5'h14 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_20_io_i_write_slot_T_2 = 5'h14 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_20_io_i_write_slot_T_5 = 5'h14 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_21_io_i_write_slot_T = 5'h15 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_21_io_i_write_slot_T_2 = 5'h15 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_21_io_i_write_slot_T_5 = 5'h15 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_22_io_i_write_slot_T = 5'h16 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_22_io_i_write_slot_T_2 = 5'h16 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_22_io_i_write_slot_T_5 = 5'h16 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_23_io_i_write_slot_T = 5'h17 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_23_io_i_write_slot_T_2 = 5'h17 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_23_io_i_write_slot_T_5 = 5'h17 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_24_io_i_write_slot_T = 5'h18 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_24_io_i_write_slot_T_2 = 5'h18 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_24_io_i_write_slot_T_5 = 5'h18 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_25_io_i_write_slot_T = 5'h19 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_25_io_i_write_slot_T_2 = 5'h19 == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_25_io_i_write_slot_T_5 = 5'h19 == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_26_io_i_write_slot_T = 5'h1a == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_26_io_i_write_slot_T_2 = 5'h1a == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_26_io_i_write_slot_T_5 = 5'h1a == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_27_io_i_write_slot_T = 5'h1b == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_27_io_i_write_slot_T_2 = 5'h1b == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_27_io_i_write_slot_T_5 = 5'h1b == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_28_io_i_write_slot_T = 5'h1c == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_28_io_i_write_slot_T_2 = 5'h1c == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_28_io_i_write_slot_T_5 = 5'h1c == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_29_io_i_write_slot_T = 5'h1d == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_29_io_i_write_slot_T_2 = 5'h1d == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_29_io_i_write_slot_T_5 = 5'h1d == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_30_io_i_write_slot_T = 5'h1e == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_30_io_i_write_slot_T_2 = 5'h1e == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_30_io_i_write_slot_T_5 = 5'h1e == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_31_io_i_write_slot_T = 5'h1f == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_31_io_i_write_slot_T_2 = 5'h1f == write_idx1 & write_idx1 != 5'h1f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_31_io_i_write_slot_T_5 = 5'h1f == write_idx2 & write_idx2 != 5'h1f; // @[reservation_station.scala 119:29]
  Reservation_Station_Slot reservation_station_0 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_0_clock),
    .reset(reservation_station_0_reset),
    .io_o_valid(reservation_station_0_io_o_valid),
    .io_o_ready_to_issue(reservation_station_0_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_0_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_0_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_0_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_0_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_0_io_i_exception),
    .io_i_write_slot(reservation_station_0_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_0_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_0_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_0_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_0_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_0_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_0_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_0_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_0_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_0_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_0_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_0_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_0_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_0_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_0_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_0_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_0_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_0_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_0_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_0_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_0_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_0_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_0_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_0_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_0_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_0_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_0_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_0_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_0_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_0_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_0_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_0_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_0_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_0_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_0_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_0_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_0_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_0_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_0_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_0_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_0_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_0_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_0_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_0_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_0_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_0_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_0_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_0_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_0_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_0_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_0_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_0_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_0_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_0_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_0_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_0_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_0_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_0_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_0_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_0_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_0_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_0_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_0_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_0_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_1 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_1_clock),
    .reset(reservation_station_1_reset),
    .io_o_valid(reservation_station_1_io_o_valid),
    .io_o_ready_to_issue(reservation_station_1_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_1_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_1_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_1_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_1_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_1_io_i_exception),
    .io_i_write_slot(reservation_station_1_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_1_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_1_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_1_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_1_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_1_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_1_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_1_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_1_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_1_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_1_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_1_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_1_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_1_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_1_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_1_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_1_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_1_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_1_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_1_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_1_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_1_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_1_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_1_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_1_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_1_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_1_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_1_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_1_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_1_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_1_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_1_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_1_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_1_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_1_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_1_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_1_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_1_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_1_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_1_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_1_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_1_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_1_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_1_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_1_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_1_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_1_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_1_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_1_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_1_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_1_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_1_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_1_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_1_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_1_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_1_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_1_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_1_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_1_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_1_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_1_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_1_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_1_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_1_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_2 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_2_clock),
    .reset(reservation_station_2_reset),
    .io_o_valid(reservation_station_2_io_o_valid),
    .io_o_ready_to_issue(reservation_station_2_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_2_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_2_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_2_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_2_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_2_io_i_exception),
    .io_i_write_slot(reservation_station_2_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_2_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_2_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_2_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_2_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_2_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_2_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_2_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_2_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_2_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_2_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_2_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_2_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_2_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_2_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_2_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_2_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_2_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_2_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_2_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_2_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_2_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_2_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_2_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_2_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_2_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_2_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_2_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_2_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_2_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_2_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_2_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_2_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_2_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_2_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_2_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_2_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_2_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_2_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_2_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_2_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_2_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_2_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_2_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_2_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_2_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_2_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_2_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_2_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_2_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_2_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_2_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_2_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_2_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_2_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_2_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_2_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_2_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_2_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_2_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_2_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_2_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_2_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_2_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_3 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_3_clock),
    .reset(reservation_station_3_reset),
    .io_o_valid(reservation_station_3_io_o_valid),
    .io_o_ready_to_issue(reservation_station_3_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_3_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_3_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_3_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_3_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_3_io_i_exception),
    .io_i_write_slot(reservation_station_3_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_3_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_3_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_3_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_3_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_3_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_3_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_3_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_3_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_3_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_3_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_3_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_3_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_3_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_3_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_3_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_3_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_3_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_3_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_3_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_3_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_3_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_3_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_3_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_3_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_3_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_3_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_3_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_3_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_3_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_3_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_3_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_3_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_3_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_3_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_3_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_3_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_3_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_3_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_3_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_3_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_3_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_3_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_3_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_3_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_3_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_3_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_3_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_3_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_3_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_3_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_3_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_3_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_3_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_3_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_3_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_3_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_3_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_3_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_3_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_3_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_3_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_3_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_3_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_4 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_4_clock),
    .reset(reservation_station_4_reset),
    .io_o_valid(reservation_station_4_io_o_valid),
    .io_o_ready_to_issue(reservation_station_4_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_4_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_4_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_4_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_4_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_4_io_i_exception),
    .io_i_write_slot(reservation_station_4_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_4_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_4_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_4_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_4_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_4_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_4_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_4_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_4_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_4_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_4_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_4_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_4_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_4_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_4_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_4_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_4_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_4_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_4_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_4_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_4_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_4_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_4_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_4_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_4_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_4_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_4_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_4_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_4_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_4_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_4_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_4_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_4_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_4_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_4_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_4_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_4_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_4_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_4_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_4_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_4_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_4_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_4_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_4_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_4_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_4_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_4_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_4_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_4_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_4_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_4_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_4_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_4_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_4_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_4_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_4_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_4_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_4_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_4_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_4_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_4_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_4_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_4_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_4_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_5 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_5_clock),
    .reset(reservation_station_5_reset),
    .io_o_valid(reservation_station_5_io_o_valid),
    .io_o_ready_to_issue(reservation_station_5_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_5_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_5_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_5_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_5_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_5_io_i_exception),
    .io_i_write_slot(reservation_station_5_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_5_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_5_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_5_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_5_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_5_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_5_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_5_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_5_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_5_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_5_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_5_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_5_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_5_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_5_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_5_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_5_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_5_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_5_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_5_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_5_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_5_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_5_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_5_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_5_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_5_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_5_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_5_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_5_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_5_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_5_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_5_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_5_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_5_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_5_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_5_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_5_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_5_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_5_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_5_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_5_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_5_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_5_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_5_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_5_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_5_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_5_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_5_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_5_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_5_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_5_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_5_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_5_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_5_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_5_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_5_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_5_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_5_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_5_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_5_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_5_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_5_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_5_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_5_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_6 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_6_clock),
    .reset(reservation_station_6_reset),
    .io_o_valid(reservation_station_6_io_o_valid),
    .io_o_ready_to_issue(reservation_station_6_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_6_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_6_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_6_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_6_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_6_io_i_exception),
    .io_i_write_slot(reservation_station_6_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_6_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_6_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_6_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_6_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_6_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_6_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_6_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_6_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_6_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_6_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_6_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_6_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_6_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_6_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_6_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_6_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_6_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_6_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_6_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_6_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_6_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_6_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_6_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_6_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_6_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_6_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_6_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_6_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_6_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_6_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_6_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_6_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_6_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_6_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_6_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_6_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_6_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_6_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_6_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_6_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_6_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_6_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_6_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_6_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_6_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_6_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_6_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_6_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_6_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_6_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_6_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_6_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_6_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_6_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_6_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_6_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_6_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_6_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_6_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_6_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_6_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_6_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_6_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_7 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_7_clock),
    .reset(reservation_station_7_reset),
    .io_o_valid(reservation_station_7_io_o_valid),
    .io_o_ready_to_issue(reservation_station_7_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_7_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_7_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_7_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_7_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_7_io_i_exception),
    .io_i_write_slot(reservation_station_7_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_7_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_7_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_7_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_7_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_7_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_7_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_7_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_7_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_7_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_7_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_7_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_7_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_7_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_7_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_7_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_7_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_7_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_7_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_7_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_7_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_7_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_7_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_7_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_7_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_7_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_7_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_7_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_7_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_7_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_7_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_7_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_7_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_7_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_7_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_7_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_7_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_7_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_7_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_7_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_7_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_7_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_7_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_7_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_7_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_7_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_7_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_7_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_7_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_7_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_7_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_7_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_7_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_7_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_7_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_7_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_7_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_7_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_7_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_7_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_7_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_7_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_7_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_7_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_8 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_8_clock),
    .reset(reservation_station_8_reset),
    .io_o_valid(reservation_station_8_io_o_valid),
    .io_o_ready_to_issue(reservation_station_8_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_8_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_8_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_8_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_8_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_8_io_i_exception),
    .io_i_write_slot(reservation_station_8_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_8_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_8_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_8_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_8_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_8_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_8_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_8_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_8_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_8_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_8_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_8_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_8_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_8_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_8_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_8_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_8_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_8_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_8_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_8_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_8_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_8_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_8_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_8_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_8_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_8_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_8_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_8_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_8_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_8_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_8_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_8_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_8_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_8_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_8_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_8_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_8_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_8_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_8_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_8_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_8_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_8_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_8_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_8_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_8_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_8_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_8_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_8_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_8_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_8_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_8_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_8_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_8_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_8_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_8_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_8_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_8_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_8_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_8_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_8_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_8_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_8_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_8_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_8_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_9 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_9_clock),
    .reset(reservation_station_9_reset),
    .io_o_valid(reservation_station_9_io_o_valid),
    .io_o_ready_to_issue(reservation_station_9_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_9_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_9_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_9_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_9_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_9_io_i_exception),
    .io_i_write_slot(reservation_station_9_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_9_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_9_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_9_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_9_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_9_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_9_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_9_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_9_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_9_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_9_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_9_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_9_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_9_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_9_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_9_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_9_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_9_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_9_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_9_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_9_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_9_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_9_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_9_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_9_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_9_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_9_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_9_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_9_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_9_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_9_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_9_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_9_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_9_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_9_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_9_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_9_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_9_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_9_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_9_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_9_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_9_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_9_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_9_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_9_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_9_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_9_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_9_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_9_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_9_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_9_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_9_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_9_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_9_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_9_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_9_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_9_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_9_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_9_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_9_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_9_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_9_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_9_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_9_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_10 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_10_clock),
    .reset(reservation_station_10_reset),
    .io_o_valid(reservation_station_10_io_o_valid),
    .io_o_ready_to_issue(reservation_station_10_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_10_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_10_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_10_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_10_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_10_io_i_exception),
    .io_i_write_slot(reservation_station_10_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_10_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_10_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_10_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_10_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_10_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_10_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_10_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_10_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_10_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_10_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_10_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_10_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_10_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_10_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_10_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_10_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_10_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_10_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_10_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_10_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_10_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_10_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_10_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_10_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_10_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_10_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_10_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_10_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_10_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_10_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_10_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_10_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_10_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_10_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_10_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_10_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_10_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_10_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_10_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_10_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_10_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_10_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_10_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_10_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_10_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_10_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_10_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_10_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_10_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_10_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_10_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_10_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_10_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_10_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_10_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_10_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_10_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_10_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_10_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_10_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_10_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_10_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_10_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_11 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_11_clock),
    .reset(reservation_station_11_reset),
    .io_o_valid(reservation_station_11_io_o_valid),
    .io_o_ready_to_issue(reservation_station_11_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_11_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_11_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_11_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_11_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_11_io_i_exception),
    .io_i_write_slot(reservation_station_11_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_11_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_11_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_11_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_11_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_11_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_11_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_11_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_11_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_11_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_11_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_11_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_11_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_11_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_11_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_11_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_11_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_11_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_11_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_11_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_11_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_11_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_11_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_11_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_11_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_11_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_11_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_11_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_11_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_11_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_11_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_11_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_11_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_11_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_11_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_11_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_11_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_11_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_11_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_11_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_11_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_11_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_11_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_11_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_11_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_11_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_11_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_11_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_11_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_11_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_11_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_11_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_11_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_11_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_11_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_11_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_11_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_11_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_11_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_11_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_11_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_11_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_11_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_11_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_12 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_12_clock),
    .reset(reservation_station_12_reset),
    .io_o_valid(reservation_station_12_io_o_valid),
    .io_o_ready_to_issue(reservation_station_12_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_12_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_12_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_12_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_12_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_12_io_i_exception),
    .io_i_write_slot(reservation_station_12_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_12_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_12_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_12_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_12_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_12_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_12_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_12_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_12_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_12_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_12_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_12_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_12_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_12_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_12_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_12_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_12_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_12_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_12_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_12_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_12_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_12_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_12_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_12_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_12_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_12_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_12_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_12_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_12_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_12_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_12_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_12_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_12_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_12_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_12_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_12_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_12_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_12_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_12_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_12_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_12_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_12_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_12_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_12_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_12_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_12_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_12_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_12_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_12_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_12_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_12_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_12_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_12_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_12_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_12_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_12_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_12_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_12_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_12_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_12_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_12_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_12_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_12_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_12_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_13 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_13_clock),
    .reset(reservation_station_13_reset),
    .io_o_valid(reservation_station_13_io_o_valid),
    .io_o_ready_to_issue(reservation_station_13_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_13_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_13_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_13_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_13_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_13_io_i_exception),
    .io_i_write_slot(reservation_station_13_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_13_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_13_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_13_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_13_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_13_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_13_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_13_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_13_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_13_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_13_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_13_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_13_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_13_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_13_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_13_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_13_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_13_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_13_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_13_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_13_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_13_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_13_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_13_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_13_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_13_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_13_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_13_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_13_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_13_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_13_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_13_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_13_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_13_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_13_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_13_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_13_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_13_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_13_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_13_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_13_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_13_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_13_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_13_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_13_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_13_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_13_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_13_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_13_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_13_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_13_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_13_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_13_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_13_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_13_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_13_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_13_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_13_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_13_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_13_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_13_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_13_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_13_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_13_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_14 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_14_clock),
    .reset(reservation_station_14_reset),
    .io_o_valid(reservation_station_14_io_o_valid),
    .io_o_ready_to_issue(reservation_station_14_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_14_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_14_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_14_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_14_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_14_io_i_exception),
    .io_i_write_slot(reservation_station_14_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_14_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_14_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_14_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_14_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_14_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_14_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_14_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_14_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_14_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_14_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_14_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_14_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_14_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_14_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_14_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_14_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_14_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_14_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_14_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_14_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_14_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_14_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_14_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_14_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_14_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_14_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_14_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_14_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_14_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_14_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_14_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_14_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_14_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_14_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_14_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_14_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_14_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_14_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_14_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_14_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_14_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_14_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_14_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_14_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_14_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_14_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_14_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_14_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_14_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_14_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_14_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_14_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_14_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_14_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_14_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_14_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_14_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_14_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_14_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_14_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_14_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_14_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_14_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_15 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_15_clock),
    .reset(reservation_station_15_reset),
    .io_o_valid(reservation_station_15_io_o_valid),
    .io_o_ready_to_issue(reservation_station_15_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_15_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_15_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_15_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_15_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_15_io_i_exception),
    .io_i_write_slot(reservation_station_15_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_15_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_15_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_15_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_15_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_15_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_15_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_15_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_15_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_15_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_15_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_15_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_15_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_15_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_15_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_15_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_15_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_15_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_15_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_15_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_15_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_15_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_15_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_15_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_15_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_15_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_15_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_15_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_15_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_15_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_15_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_15_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_15_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_15_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_15_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_15_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_15_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_15_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_15_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_15_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_15_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_15_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_15_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_15_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_15_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_15_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_15_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_15_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_15_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_15_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_15_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_15_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_15_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_15_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_15_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_15_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_15_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_15_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_15_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_15_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_15_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_15_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_15_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_15_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_16 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_16_clock),
    .reset(reservation_station_16_reset),
    .io_o_valid(reservation_station_16_io_o_valid),
    .io_o_ready_to_issue(reservation_station_16_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_16_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_16_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_16_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_16_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_16_io_i_exception),
    .io_i_write_slot(reservation_station_16_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_16_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_16_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_16_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_16_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_16_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_16_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_16_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_16_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_16_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_16_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_16_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_16_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_16_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_16_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_16_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_16_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_16_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_16_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_16_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_16_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_16_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_16_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_16_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_16_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_16_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_16_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_16_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_16_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_16_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_16_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_16_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_16_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_16_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_16_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_16_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_16_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_16_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_16_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_16_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_16_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_16_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_16_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_16_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_16_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_16_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_16_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_16_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_16_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_16_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_16_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_16_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_16_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_16_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_16_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_16_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_16_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_16_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_16_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_16_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_16_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_16_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_16_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_16_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_17 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_17_clock),
    .reset(reservation_station_17_reset),
    .io_o_valid(reservation_station_17_io_o_valid),
    .io_o_ready_to_issue(reservation_station_17_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_17_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_17_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_17_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_17_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_17_io_i_exception),
    .io_i_write_slot(reservation_station_17_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_17_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_17_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_17_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_17_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_17_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_17_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_17_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_17_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_17_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_17_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_17_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_17_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_17_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_17_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_17_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_17_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_17_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_17_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_17_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_17_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_17_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_17_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_17_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_17_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_17_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_17_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_17_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_17_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_17_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_17_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_17_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_17_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_17_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_17_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_17_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_17_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_17_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_17_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_17_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_17_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_17_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_17_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_17_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_17_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_17_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_17_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_17_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_17_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_17_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_17_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_17_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_17_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_17_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_17_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_17_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_17_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_17_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_17_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_17_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_17_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_17_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_17_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_17_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_18 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_18_clock),
    .reset(reservation_station_18_reset),
    .io_o_valid(reservation_station_18_io_o_valid),
    .io_o_ready_to_issue(reservation_station_18_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_18_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_18_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_18_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_18_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_18_io_i_exception),
    .io_i_write_slot(reservation_station_18_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_18_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_18_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_18_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_18_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_18_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_18_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_18_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_18_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_18_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_18_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_18_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_18_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_18_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_18_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_18_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_18_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_18_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_18_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_18_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_18_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_18_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_18_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_18_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_18_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_18_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_18_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_18_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_18_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_18_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_18_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_18_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_18_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_18_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_18_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_18_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_18_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_18_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_18_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_18_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_18_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_18_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_18_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_18_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_18_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_18_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_18_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_18_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_18_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_18_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_18_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_18_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_18_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_18_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_18_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_18_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_18_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_18_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_18_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_18_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_18_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_18_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_18_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_18_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_19 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_19_clock),
    .reset(reservation_station_19_reset),
    .io_o_valid(reservation_station_19_io_o_valid),
    .io_o_ready_to_issue(reservation_station_19_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_19_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_19_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_19_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_19_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_19_io_i_exception),
    .io_i_write_slot(reservation_station_19_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_19_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_19_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_19_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_19_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_19_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_19_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_19_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_19_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_19_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_19_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_19_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_19_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_19_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_19_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_19_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_19_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_19_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_19_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_19_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_19_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_19_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_19_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_19_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_19_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_19_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_19_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_19_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_19_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_19_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_19_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_19_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_19_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_19_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_19_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_19_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_19_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_19_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_19_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_19_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_19_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_19_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_19_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_19_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_19_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_19_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_19_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_19_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_19_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_19_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_19_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_19_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_19_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_19_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_19_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_19_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_19_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_19_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_19_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_19_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_19_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_19_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_19_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_19_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_20 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_20_clock),
    .reset(reservation_station_20_reset),
    .io_o_valid(reservation_station_20_io_o_valid),
    .io_o_ready_to_issue(reservation_station_20_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_20_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_20_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_20_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_20_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_20_io_i_exception),
    .io_i_write_slot(reservation_station_20_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_20_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_20_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_20_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_20_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_20_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_20_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_20_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_20_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_20_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_20_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_20_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_20_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_20_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_20_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_20_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_20_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_20_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_20_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_20_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_20_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_20_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_20_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_20_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_20_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_20_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_20_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_20_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_20_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_20_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_20_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_20_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_20_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_20_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_20_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_20_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_20_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_20_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_20_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_20_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_20_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_20_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_20_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_20_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_20_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_20_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_20_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_20_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_20_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_20_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_20_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_20_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_20_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_20_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_20_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_20_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_20_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_20_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_20_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_20_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_20_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_20_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_20_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_20_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_21 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_21_clock),
    .reset(reservation_station_21_reset),
    .io_o_valid(reservation_station_21_io_o_valid),
    .io_o_ready_to_issue(reservation_station_21_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_21_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_21_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_21_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_21_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_21_io_i_exception),
    .io_i_write_slot(reservation_station_21_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_21_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_21_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_21_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_21_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_21_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_21_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_21_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_21_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_21_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_21_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_21_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_21_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_21_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_21_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_21_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_21_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_21_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_21_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_21_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_21_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_21_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_21_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_21_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_21_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_21_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_21_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_21_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_21_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_21_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_21_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_21_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_21_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_21_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_21_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_21_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_21_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_21_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_21_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_21_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_21_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_21_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_21_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_21_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_21_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_21_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_21_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_21_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_21_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_21_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_21_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_21_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_21_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_21_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_21_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_21_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_21_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_21_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_21_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_21_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_21_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_21_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_21_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_21_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_22 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_22_clock),
    .reset(reservation_station_22_reset),
    .io_o_valid(reservation_station_22_io_o_valid),
    .io_o_ready_to_issue(reservation_station_22_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_22_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_22_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_22_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_22_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_22_io_i_exception),
    .io_i_write_slot(reservation_station_22_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_22_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_22_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_22_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_22_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_22_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_22_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_22_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_22_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_22_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_22_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_22_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_22_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_22_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_22_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_22_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_22_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_22_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_22_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_22_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_22_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_22_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_22_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_22_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_22_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_22_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_22_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_22_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_22_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_22_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_22_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_22_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_22_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_22_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_22_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_22_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_22_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_22_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_22_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_22_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_22_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_22_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_22_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_22_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_22_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_22_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_22_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_22_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_22_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_22_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_22_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_22_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_22_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_22_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_22_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_22_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_22_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_22_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_22_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_22_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_22_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_22_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_22_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_22_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_23 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_23_clock),
    .reset(reservation_station_23_reset),
    .io_o_valid(reservation_station_23_io_o_valid),
    .io_o_ready_to_issue(reservation_station_23_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_23_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_23_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_23_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_23_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_23_io_i_exception),
    .io_i_write_slot(reservation_station_23_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_23_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_23_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_23_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_23_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_23_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_23_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_23_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_23_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_23_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_23_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_23_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_23_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_23_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_23_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_23_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_23_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_23_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_23_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_23_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_23_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_23_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_23_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_23_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_23_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_23_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_23_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_23_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_23_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_23_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_23_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_23_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_23_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_23_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_23_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_23_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_23_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_23_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_23_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_23_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_23_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_23_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_23_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_23_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_23_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_23_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_23_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_23_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_23_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_23_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_23_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_23_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_23_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_23_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_23_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_23_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_23_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_23_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_23_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_23_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_23_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_23_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_23_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_23_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_24 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_24_clock),
    .reset(reservation_station_24_reset),
    .io_o_valid(reservation_station_24_io_o_valid),
    .io_o_ready_to_issue(reservation_station_24_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_24_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_24_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_24_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_24_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_24_io_i_exception),
    .io_i_write_slot(reservation_station_24_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_24_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_24_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_24_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_24_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_24_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_24_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_24_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_24_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_24_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_24_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_24_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_24_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_24_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_24_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_24_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_24_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_24_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_24_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_24_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_24_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_24_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_24_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_24_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_24_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_24_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_24_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_24_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_24_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_24_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_24_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_24_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_24_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_24_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_24_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_24_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_24_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_24_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_24_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_24_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_24_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_24_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_24_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_24_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_24_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_24_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_24_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_24_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_24_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_24_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_24_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_24_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_24_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_24_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_24_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_24_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_24_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_24_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_24_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_24_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_24_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_24_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_24_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_24_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_25 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_25_clock),
    .reset(reservation_station_25_reset),
    .io_o_valid(reservation_station_25_io_o_valid),
    .io_o_ready_to_issue(reservation_station_25_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_25_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_25_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_25_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_25_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_25_io_i_exception),
    .io_i_write_slot(reservation_station_25_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_25_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_25_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_25_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_25_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_25_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_25_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_25_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_25_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_25_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_25_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_25_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_25_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_25_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_25_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_25_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_25_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_25_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_25_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_25_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_25_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_25_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_25_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_25_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_25_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_25_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_25_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_25_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_25_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_25_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_25_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_25_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_25_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_25_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_25_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_25_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_25_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_25_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_25_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_25_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_25_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_25_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_25_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_25_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_25_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_25_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_25_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_25_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_25_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_25_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_25_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_25_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_25_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_25_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_25_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_25_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_25_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_25_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_25_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_25_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_25_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_25_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_25_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_25_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_26 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_26_clock),
    .reset(reservation_station_26_reset),
    .io_o_valid(reservation_station_26_io_o_valid),
    .io_o_ready_to_issue(reservation_station_26_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_26_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_26_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_26_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_26_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_26_io_i_exception),
    .io_i_write_slot(reservation_station_26_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_26_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_26_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_26_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_26_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_26_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_26_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_26_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_26_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_26_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_26_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_26_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_26_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_26_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_26_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_26_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_26_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_26_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_26_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_26_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_26_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_26_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_26_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_26_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_26_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_26_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_26_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_26_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_26_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_26_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_26_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_26_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_26_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_26_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_26_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_26_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_26_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_26_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_26_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_26_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_26_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_26_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_26_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_26_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_26_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_26_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_26_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_26_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_26_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_26_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_26_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_26_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_26_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_26_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_26_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_26_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_26_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_26_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_26_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_26_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_26_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_26_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_26_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_26_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_27 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_27_clock),
    .reset(reservation_station_27_reset),
    .io_o_valid(reservation_station_27_io_o_valid),
    .io_o_ready_to_issue(reservation_station_27_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_27_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_27_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_27_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_27_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_27_io_i_exception),
    .io_i_write_slot(reservation_station_27_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_27_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_27_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_27_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_27_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_27_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_27_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_27_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_27_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_27_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_27_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_27_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_27_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_27_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_27_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_27_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_27_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_27_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_27_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_27_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_27_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_27_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_27_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_27_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_27_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_27_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_27_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_27_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_27_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_27_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_27_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_27_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_27_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_27_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_27_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_27_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_27_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_27_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_27_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_27_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_27_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_27_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_27_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_27_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_27_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_27_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_27_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_27_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_27_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_27_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_27_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_27_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_27_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_27_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_27_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_27_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_27_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_27_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_27_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_27_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_27_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_27_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_27_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_27_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_28 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_28_clock),
    .reset(reservation_station_28_reset),
    .io_o_valid(reservation_station_28_io_o_valid),
    .io_o_ready_to_issue(reservation_station_28_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_28_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_28_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_28_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_28_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_28_io_i_exception),
    .io_i_write_slot(reservation_station_28_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_28_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_28_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_28_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_28_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_28_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_28_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_28_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_28_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_28_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_28_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_28_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_28_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_28_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_28_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_28_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_28_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_28_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_28_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_28_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_28_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_28_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_28_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_28_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_28_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_28_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_28_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_28_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_28_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_28_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_28_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_28_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_28_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_28_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_28_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_28_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_28_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_28_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_28_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_28_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_28_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_28_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_28_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_28_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_28_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_28_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_28_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_28_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_28_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_28_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_28_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_28_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_28_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_28_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_28_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_28_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_28_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_28_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_28_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_28_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_28_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_28_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_28_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_28_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_29 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_29_clock),
    .reset(reservation_station_29_reset),
    .io_o_valid(reservation_station_29_io_o_valid),
    .io_o_ready_to_issue(reservation_station_29_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_29_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_29_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_29_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_29_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_29_io_i_exception),
    .io_i_write_slot(reservation_station_29_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_29_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_29_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_29_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_29_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_29_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_29_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_29_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_29_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_29_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_29_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_29_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_29_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_29_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_29_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_29_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_29_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_29_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_29_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_29_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_29_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_29_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_29_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_29_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_29_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_29_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_29_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_29_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_29_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_29_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_29_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_29_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_29_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_29_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_29_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_29_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_29_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_29_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_29_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_29_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_29_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_29_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_29_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_29_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_29_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_29_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_29_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_29_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_29_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_29_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_29_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_29_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_29_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_29_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_29_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_29_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_29_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_29_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_29_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_29_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_29_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_29_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_29_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_29_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_30 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_30_clock),
    .reset(reservation_station_30_reset),
    .io_o_valid(reservation_station_30_io_o_valid),
    .io_o_ready_to_issue(reservation_station_30_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_30_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_30_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_30_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_30_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_30_io_i_exception),
    .io_i_write_slot(reservation_station_30_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_30_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_30_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_30_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_30_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_30_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_30_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_30_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_30_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_30_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_30_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_30_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_30_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_30_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_30_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_30_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_30_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_30_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_30_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_30_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_30_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_30_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_30_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_30_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_30_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_30_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_30_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_30_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_30_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_30_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_30_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_30_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_30_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_30_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_30_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_30_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_30_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_30_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_30_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_30_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_30_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_30_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_30_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_30_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_30_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_30_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_30_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_30_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_30_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_30_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_30_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_30_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_30_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_30_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_30_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_30_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_30_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_30_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_30_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_30_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_30_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_30_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_30_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_30_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_31 ( // @[reservation_station.scala 38:56]
    .clock(reservation_station_31_clock),
    .reset(reservation_station_31_reset),
    .io_o_valid(reservation_station_31_io_o_valid),
    .io_o_ready_to_issue(reservation_station_31_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_31_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_31_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_31_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_31_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_31_io_i_exception),
    .io_i_write_slot(reservation_station_31_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_31_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_31_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_31_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_31_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_31_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_31_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_31_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_31_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_31_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_31_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_31_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_31_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_31_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_31_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_31_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_31_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_31_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_31_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_31_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_31_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_31_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_31_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_31_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_31_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_31_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_31_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_31_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_31_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_31_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_31_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_31_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_31_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_31_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_31_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_31_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_31_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_31_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_31_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_31_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_31_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_31_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_31_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_31_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_31_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_31_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_31_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_31_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_31_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_31_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_31_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_31_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_31_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_31_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_31_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_31_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_31_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_31_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_31_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_31_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_31_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_31_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_31_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_31_io_i_ROB_first_entry)
  );
  assign io_o_issue_packs_0_valid = issue_num == 2'h1 | issue_num == 2'h2; // @[reservation_station.scala 93:38]
  assign io_o_issue_packs_0_pc = _issue1_func_code_T ? reservation_station_0_io_o_uop_pc : _io_o_issue_packs_0_T_62_pc; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_inst = _issue1_func_code_T ? reservation_station_0_io_o_uop_inst :
    _io_o_issue_packs_0_T_62_inst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_func_code = _issue1_func_code_T ? reservation_station_0_io_o_uop_func_code :
    _io_o_issue_packs_0_T_62_func_code; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_valid = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_62_branch_predict_pack_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_target = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_62_branch_predict_pack_target; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_branch_type = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_62_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_select = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_62_branch_predict_pack_select; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_taken = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_62_branch_predict_pack_taken; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_62_phy_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_stale_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_62_stale_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_62_arch_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_inst_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_62_inst_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_regWen = _issue1_func_code_T ? reservation_station_0_io_o_uop_regWen :
    _io_o_issue_packs_0_T_62_regWen; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src1_valid = _issue1_func_code_T ? reservation_station_0_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_62_src1_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_rs1 = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_62_phy_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_rs1 = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_62_arch_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src2_valid = _issue1_func_code_T ? reservation_station_0_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_62_src2_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_rs2 = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_62_phy_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_rs2 = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_62_arch_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_rob_idx = _issue1_func_code_T ? reservation_station_0_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_62_rob_idx; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_imm = _issue1_func_code_T ? reservation_station_0_io_o_uop_imm :
    _io_o_issue_packs_0_T_62_imm; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src1_value = _issue1_func_code_T ? reservation_station_0_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_62_src1_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src2_value = _issue1_func_code_T ? reservation_station_0_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_62_src2_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_op1_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_62_op1_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_op2_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_62_op2_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_alu_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_62_alu_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_branch_type :
    _io_o_issue_packs_0_T_62_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_mem_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_62_mem_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_valid = issue_num == 2'h2; // @[reservation_station.scala 94:31]
  assign io_o_issue_packs_1_pc = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_pc : _io_o_issue_packs_1_T_62_pc
    ; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_inst = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_inst :
    _io_o_issue_packs_1_T_62_inst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_func_code = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_func_code :
    _io_o_issue_packs_1_T_62_func_code; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_valid = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_62_branch_predict_pack_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_target = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_62_branch_predict_pack_target; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_branch_type = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_62_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_select = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_62_branch_predict_pack_select; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_taken = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_62_branch_predict_pack_taken; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_dst = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_62_phy_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_stale_dst = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_62_stale_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_dst = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_62_arch_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_inst_type = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_62_inst_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_regWen = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_regWen :
    _io_o_issue_packs_1_T_62_regWen; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src1_valid = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_62_src1_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_rs1 = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_62_phy_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_rs1 = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_62_arch_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src2_valid = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_62_src2_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_rs2 = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_62_phy_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_rs2 = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_62_arch_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_rob_idx = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_62_rob_idx; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_imm = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_imm :
    _io_o_issue_packs_1_T_62_imm; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src1_value = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_src1_value :
    _io_o_issue_packs_1_T_62_src1_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src2_value = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_src2_value :
    _io_o_issue_packs_1_T_62_src2_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_op1_sel = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_62_op1_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_op2_sel = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_62_op2_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_alu_sel = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_62_alu_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_type = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_branch_type :
    _io_o_issue_packs_1_T_62_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_mem_type = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_62_mem_type; // @[Mux.scala 101:16]
  assign io_o_full = _write_num_T | _write_num_T_1; // @[reservation_station.scala 104:47]
  assign reservation_station_0_clock = clock;
  assign reservation_station_0_reset = reset;
  assign reservation_station_0_io_i_issue_granted = (_issue1_func_code_T | _io_o_issue_packs_1_T) & ~(io_i_exception |
    io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_0_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_0_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_0_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_0_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_0_io_i_write_slot = _reservation_station_0_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_0_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_0_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_0_io_i_uop_valid = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_pc = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_inst = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_func_code = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_target = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_branch_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_select = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_taken = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_phy_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_stale_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_arch_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_inst_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_regWen = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_src1_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_phy_rs1 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_arch_rs1 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_src2_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_phy_rs2 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_arch_rs2 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_rob_idx = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_imm = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_src1_value = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_src2_value = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_op1_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_op2_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_alu_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_mem_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_0_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_0_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_0_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_0_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_1_clock = clock;
  assign reservation_station_1_reset = reset;
  assign reservation_station_1_io_i_issue_granted = (_issue1_func_code_T_1 | _io_o_issue_packs_1_T_1) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_1_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_1_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_1_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_1_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_1_io_i_write_slot = _reservation_station_1_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_1_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_1_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_1_io_i_uop_valid = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_pc = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_inst = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_func_code = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_target = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_branch_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_select = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_taken = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_phy_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_stale_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_arch_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_inst_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_regWen = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_src1_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_phy_rs1 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_arch_rs1 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_src2_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_phy_rs2 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_arch_rs2 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_rob_idx = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_imm = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_src1_value = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_src2_value = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_op1_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_op2_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_alu_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_mem_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_1_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_1_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_1_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_1_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_2_clock = clock;
  assign reservation_station_2_reset = reset;
  assign reservation_station_2_io_i_issue_granted = (_issue1_func_code_T_2 | _io_o_issue_packs_1_T_2) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_2_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_2_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_2_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_2_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_2_io_i_write_slot = _reservation_station_2_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_2_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_2_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_2_io_i_uop_valid = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_pc = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_inst = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_func_code = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_target = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_branch_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_select = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_taken = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_phy_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_stale_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_arch_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_inst_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_regWen = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_src1_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_phy_rs1 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_arch_rs1 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_src2_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_phy_rs2 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_arch_rs2 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_rob_idx = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_imm = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_src1_value = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_src2_value = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_op1_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_op2_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_alu_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_mem_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_2_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_2_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_2_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_2_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_3_clock = clock;
  assign reservation_station_3_reset = reset;
  assign reservation_station_3_io_i_issue_granted = (_issue1_func_code_T_3 | _io_o_issue_packs_1_T_3) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_3_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_3_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_3_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_3_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_3_io_i_write_slot = _reservation_station_3_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_3_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_3_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_3_io_i_uop_valid = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_pc = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_inst = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_func_code = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_target = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_branch_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_select = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_taken = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_phy_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_stale_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_arch_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_inst_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_regWen = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_src1_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_phy_rs1 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_arch_rs1 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_src2_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_phy_rs2 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_arch_rs2 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_rob_idx = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_imm = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_src1_value = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_src2_value = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_op1_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_op2_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_alu_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_mem_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_3_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_3_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_3_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_3_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_4_clock = clock;
  assign reservation_station_4_reset = reset;
  assign reservation_station_4_io_i_issue_granted = (_issue1_func_code_T_4 | _io_o_issue_packs_1_T_4) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_4_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_4_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_4_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_4_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_4_io_i_write_slot = _reservation_station_4_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_4_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_4_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_4_io_i_uop_valid = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_pc = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_inst = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_func_code = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_target = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_branch_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_select = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_taken = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_phy_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_stale_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_arch_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_inst_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_regWen = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_src1_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_phy_rs1 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_arch_rs1 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_src2_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_phy_rs2 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_arch_rs2 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_rob_idx = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_imm = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_src1_value = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_src2_value = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_op1_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_op2_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_alu_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_mem_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_4_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_4_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_4_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_4_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_5_clock = clock;
  assign reservation_station_5_reset = reset;
  assign reservation_station_5_io_i_issue_granted = (_issue1_func_code_T_5 | _io_o_issue_packs_1_T_5) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_5_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_5_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_5_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_5_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_5_io_i_write_slot = _reservation_station_5_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_5_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_5_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_5_io_i_uop_valid = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_pc = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_inst = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_func_code = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_target = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_branch_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_select = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_taken = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_phy_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_stale_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_arch_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_inst_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_regWen = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_src1_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_phy_rs1 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_arch_rs1 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_src2_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_phy_rs2 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_arch_rs2 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_rob_idx = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_imm = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_src1_value = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_src2_value = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_op1_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_op2_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_alu_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_mem_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_5_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_5_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_5_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_5_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_6_clock = clock;
  assign reservation_station_6_reset = reset;
  assign reservation_station_6_io_i_issue_granted = (_issue1_func_code_T_6 | _io_o_issue_packs_1_T_6) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_6_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_6_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_6_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_6_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_6_io_i_write_slot = _reservation_station_6_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_6_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_6_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_6_io_i_uop_valid = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_pc = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_inst = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_func_code = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_target = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_branch_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_select = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_taken = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_phy_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_stale_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_arch_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_inst_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_regWen = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_src1_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_phy_rs1 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_arch_rs1 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_src2_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_phy_rs2 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_arch_rs2 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_rob_idx = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_imm = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_src1_value = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_src2_value = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_op1_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_op2_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_alu_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_mem_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_6_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_6_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_6_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_6_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_7_clock = clock;
  assign reservation_station_7_reset = reset;
  assign reservation_station_7_io_i_issue_granted = (_issue1_func_code_T_7 | _io_o_issue_packs_1_T_7) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_7_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_7_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_7_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_7_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_7_io_i_write_slot = _reservation_station_7_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_7_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_7_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_7_io_i_uop_valid = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_pc = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_inst = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_func_code = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_target = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_branch_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_select = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_taken = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_phy_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_stale_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_arch_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_inst_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_regWen = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_src1_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_phy_rs1 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_arch_rs1 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_src2_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_phy_rs2 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_arch_rs2 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_rob_idx = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_imm = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_src1_value = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_src2_value = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_op1_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_op2_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_alu_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_mem_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_7_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_7_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_7_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_7_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_8_clock = clock;
  assign reservation_station_8_reset = reset;
  assign reservation_station_8_io_i_issue_granted = (_issue1_func_code_T_8 | _io_o_issue_packs_1_T_8) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_8_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_8_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_8_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_8_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_8_io_i_write_slot = _reservation_station_8_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_8_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_8_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_8_io_i_uop_valid = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_pc = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_inst = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_func_code = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_target = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_branch_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_select = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_taken = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_phy_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_stale_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_arch_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_inst_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_regWen = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_src1_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_phy_rs1 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_arch_rs1 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_src2_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_phy_rs2 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_arch_rs2 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_rob_idx = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_imm = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_src1_value = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_src2_value = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_op1_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_op2_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_alu_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_mem_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_8_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_8_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_8_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_8_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_9_clock = clock;
  assign reservation_station_9_reset = reset;
  assign reservation_station_9_io_i_issue_granted = (_issue1_func_code_T_9 | _io_o_issue_packs_1_T_9) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_9_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_9_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_9_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_9_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_9_io_i_write_slot = _reservation_station_9_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_9_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_9_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_9_io_i_uop_valid = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_pc = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_inst = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_func_code = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_target = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_branch_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_select = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_taken = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_phy_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_stale_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_arch_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_inst_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_regWen = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_src1_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_phy_rs1 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_arch_rs1 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_src2_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_phy_rs2 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_arch_rs2 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_rob_idx = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_imm = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_src1_value = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_src2_value = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_op1_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_op2_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_alu_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_mem_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_9_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_9_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_9_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_9_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_10_clock = clock;
  assign reservation_station_10_reset = reset;
  assign reservation_station_10_io_i_issue_granted = (_issue1_func_code_T_10 | _io_o_issue_packs_1_T_10) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_10_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_10_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_10_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_10_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_10_io_i_write_slot = _reservation_station_10_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_10_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_10_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_10_io_i_uop_valid = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_pc = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_inst = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_func_code = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_target = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_branch_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_select = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_taken = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_phy_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_stale_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_arch_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_inst_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_regWen = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_src1_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_phy_rs1 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_arch_rs1 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_src2_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_phy_rs2 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_arch_rs2 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_rob_idx = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_imm = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_src1_value = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_src2_value = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_op1_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_op2_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_alu_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_mem_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_10_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_10_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_10_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_10_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_11_clock = clock;
  assign reservation_station_11_reset = reset;
  assign reservation_station_11_io_i_issue_granted = (_issue1_func_code_T_11 | _io_o_issue_packs_1_T_11) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_11_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_11_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_11_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_11_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_11_io_i_write_slot = _reservation_station_11_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_11_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_11_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_11_io_i_uop_valid = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_pc = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_inst = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_func_code = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_target = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_branch_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_select = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_taken = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_phy_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_stale_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_arch_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_inst_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_regWen = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_src1_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_phy_rs1 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_arch_rs1 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_src2_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_phy_rs2 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_arch_rs2 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_rob_idx = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_imm = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_src1_value = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_src2_value = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_op1_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_op2_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_alu_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_mem_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_11_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_11_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_11_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_11_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_12_clock = clock;
  assign reservation_station_12_reset = reset;
  assign reservation_station_12_io_i_issue_granted = (_issue1_func_code_T_12 | _io_o_issue_packs_1_T_12) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_12_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_12_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_12_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_12_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_12_io_i_write_slot = _reservation_station_12_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_12_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_12_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_12_io_i_uop_valid = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_pc = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_inst = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_func_code = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_target = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_branch_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_select = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_taken = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_phy_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_stale_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_arch_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_inst_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_regWen = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_src1_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_phy_rs1 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_arch_rs1 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_src2_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_phy_rs2 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_arch_rs2 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_rob_idx = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_imm = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_src1_value = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_src2_value = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_op1_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_op2_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_alu_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_mem_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_12_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_12_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_12_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_12_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_13_clock = clock;
  assign reservation_station_13_reset = reset;
  assign reservation_station_13_io_i_issue_granted = (_issue1_func_code_T_13 | _io_o_issue_packs_1_T_13) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_13_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_13_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_13_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_13_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_13_io_i_write_slot = _reservation_station_13_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_13_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_13_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_13_io_i_uop_valid = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_pc = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_inst = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_func_code = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_target = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_branch_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_select = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_taken = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_phy_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_stale_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_arch_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_inst_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_regWen = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_src1_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_phy_rs1 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_arch_rs1 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_src2_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_phy_rs2 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_arch_rs2 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_rob_idx = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_imm = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_src1_value = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_src2_value = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_op1_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_op2_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_alu_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_mem_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_13_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_13_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_13_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_13_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_14_clock = clock;
  assign reservation_station_14_reset = reset;
  assign reservation_station_14_io_i_issue_granted = (_issue1_func_code_T_14 | _io_o_issue_packs_1_T_14) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_14_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_14_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_14_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_14_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_14_io_i_write_slot = _reservation_station_14_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_14_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_14_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_14_io_i_uop_valid = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_pc = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_inst = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_func_code = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_target = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_branch_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_select = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_taken = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_phy_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_stale_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_arch_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_inst_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_regWen = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_src1_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_phy_rs1 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_arch_rs1 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_src2_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_phy_rs2 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_arch_rs2 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_rob_idx = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_imm = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_src1_value = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_src2_value = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_op1_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_op2_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_alu_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_mem_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_14_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_14_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_14_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_14_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_15_clock = clock;
  assign reservation_station_15_reset = reset;
  assign reservation_station_15_io_i_issue_granted = (_issue1_func_code_T_15 | _io_o_issue_packs_1_T_15) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_15_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_15_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_15_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_15_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_15_io_i_write_slot = _reservation_station_15_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_15_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_15_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_15_io_i_uop_valid = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_pc = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_inst = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_func_code = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_target = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_branch_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_select = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_taken = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_phy_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_stale_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_arch_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_inst_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_regWen = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_src1_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_phy_rs1 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_arch_rs1 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_src2_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_phy_rs2 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_arch_rs2 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_rob_idx = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_imm = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_src1_value = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_src2_value = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_op1_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_op2_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_alu_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_mem_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_15_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_15_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_15_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_15_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_16_clock = clock;
  assign reservation_station_16_reset = reset;
  assign reservation_station_16_io_i_issue_granted = (_issue1_func_code_T_16 | _io_o_issue_packs_1_T_16) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_16_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_16_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_16_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_16_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_16_io_i_write_slot = _reservation_station_16_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_16_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_16_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_16_io_i_uop_valid = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_pc = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_inst = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_func_code = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_target = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_branch_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_select = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_taken = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_phy_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_stale_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_arch_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_inst_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_regWen = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_src1_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_phy_rs1 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_arch_rs1 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_src2_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_phy_rs2 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_arch_rs2 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_rob_idx = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_imm = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_src1_value = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_src2_value = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_op1_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_op2_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_alu_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_mem_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_16_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_16_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_16_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_16_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_17_clock = clock;
  assign reservation_station_17_reset = reset;
  assign reservation_station_17_io_i_issue_granted = (_issue1_func_code_T_17 | _io_o_issue_packs_1_T_17) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_17_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_17_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_17_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_17_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_17_io_i_write_slot = _reservation_station_17_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_17_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_17_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_17_io_i_uop_valid = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_pc = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_inst = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_func_code = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_target = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_branch_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_select = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_taken = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_phy_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_stale_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_arch_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_inst_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_regWen = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_src1_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_phy_rs1 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_arch_rs1 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_src2_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_phy_rs2 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_arch_rs2 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_rob_idx = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_imm = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_src1_value = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_src2_value = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_op1_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_op2_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_alu_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_mem_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_17_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_17_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_17_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_17_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_18_clock = clock;
  assign reservation_station_18_reset = reset;
  assign reservation_station_18_io_i_issue_granted = (_issue1_func_code_T_18 | _io_o_issue_packs_1_T_18) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_18_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_18_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_18_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_18_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_18_io_i_write_slot = _reservation_station_18_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_18_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_18_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_18_io_i_uop_valid = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_pc = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_inst = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_func_code = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_target = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_branch_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_select = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_taken = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_phy_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_stale_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_arch_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_inst_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_regWen = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_src1_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_phy_rs1 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_arch_rs1 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_src2_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_phy_rs2 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_arch_rs2 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_rob_idx = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_imm = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_src1_value = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_src2_value = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_op1_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_op2_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_alu_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_mem_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_18_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_18_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_18_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_18_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_19_clock = clock;
  assign reservation_station_19_reset = reset;
  assign reservation_station_19_io_i_issue_granted = (_issue1_func_code_T_19 | _io_o_issue_packs_1_T_19) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_19_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_19_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_19_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_19_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_19_io_i_write_slot = _reservation_station_19_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_19_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_19_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_19_io_i_uop_valid = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_pc = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_inst = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_func_code = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_target = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_branch_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_select = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_taken = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_phy_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_stale_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_arch_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_inst_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_regWen = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_src1_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_phy_rs1 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_arch_rs1 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_src2_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_phy_rs2 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_arch_rs2 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_rob_idx = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_imm = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_src1_value = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_src2_value = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_op1_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_op2_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_alu_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_mem_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_19_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_19_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_19_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_19_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_20_clock = clock;
  assign reservation_station_20_reset = reset;
  assign reservation_station_20_io_i_issue_granted = (_issue1_func_code_T_20 | _io_o_issue_packs_1_T_20) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_20_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_20_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_20_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_20_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_20_io_i_write_slot = _reservation_station_20_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_20_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_20_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_20_io_i_uop_valid = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_pc = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_inst = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_func_code = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_target = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_branch_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_select = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_taken = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_phy_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_stale_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_arch_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_inst_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_regWen = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_src1_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_phy_rs1 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_arch_rs1 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_src2_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_phy_rs2 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_arch_rs2 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_rob_idx = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_imm = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_src1_value = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_src2_value = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_op1_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_op2_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_alu_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_mem_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_20_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_20_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_20_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_20_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_21_clock = clock;
  assign reservation_station_21_reset = reset;
  assign reservation_station_21_io_i_issue_granted = (_issue1_func_code_T_21 | _io_o_issue_packs_1_T_21) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_21_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_21_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_21_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_21_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_21_io_i_write_slot = _reservation_station_21_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_21_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_21_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_21_io_i_uop_valid = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_pc = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_inst = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_func_code = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_target = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_branch_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_select = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_taken = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_phy_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_stale_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_arch_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_inst_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_regWen = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_src1_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_phy_rs1 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_arch_rs1 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_src2_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_phy_rs2 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_arch_rs2 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_rob_idx = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_imm = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_src1_value = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_src2_value = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_op1_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_op2_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_alu_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_mem_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_21_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_21_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_21_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_21_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_22_clock = clock;
  assign reservation_station_22_reset = reset;
  assign reservation_station_22_io_i_issue_granted = (_issue1_func_code_T_22 | _io_o_issue_packs_1_T_22) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_22_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_22_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_22_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_22_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_22_io_i_write_slot = _reservation_station_22_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_22_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_22_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_22_io_i_uop_valid = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_pc = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_inst = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_func_code = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_target = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_branch_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_select = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_taken = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_phy_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_stale_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_arch_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_inst_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_regWen = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_src1_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_phy_rs1 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_arch_rs1 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_src2_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_phy_rs2 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_arch_rs2 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_rob_idx = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_imm = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_src1_value = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_src2_value = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_op1_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_op2_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_alu_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_mem_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_22_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_22_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_22_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_22_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_23_clock = clock;
  assign reservation_station_23_reset = reset;
  assign reservation_station_23_io_i_issue_granted = (_issue1_func_code_T_23 | _io_o_issue_packs_1_T_23) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_23_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_23_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_23_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_23_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_23_io_i_write_slot = _reservation_station_23_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_23_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_23_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_23_io_i_uop_valid = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_pc = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_inst = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_func_code = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_target = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_branch_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_select = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_taken = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_phy_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_stale_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_arch_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_inst_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_regWen = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_src1_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_phy_rs1 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_arch_rs1 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_src2_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_phy_rs2 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_arch_rs2 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_rob_idx = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_imm = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_src1_value = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_src2_value = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_op1_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_op2_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_alu_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_mem_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_23_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_23_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_23_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_23_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_24_clock = clock;
  assign reservation_station_24_reset = reset;
  assign reservation_station_24_io_i_issue_granted = (_issue1_func_code_T_24 | _io_o_issue_packs_1_T_24) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_24_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_24_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_24_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_24_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_24_io_i_write_slot = _reservation_station_24_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_24_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_24_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_24_io_i_uop_valid = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_pc = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_inst = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_func_code = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_target = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_branch_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_select = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_taken = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_phy_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_stale_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_arch_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_inst_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_regWen = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_src1_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_phy_rs1 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_arch_rs1 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_src2_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_phy_rs2 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_arch_rs2 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_rob_idx = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_imm = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_src1_value = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_src2_value = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_op1_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_op2_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_alu_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_mem_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_24_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_24_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_24_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_24_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_25_clock = clock;
  assign reservation_station_25_reset = reset;
  assign reservation_station_25_io_i_issue_granted = (_issue1_func_code_T_25 | _io_o_issue_packs_1_T_25) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_25_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_25_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_25_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_25_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_25_io_i_write_slot = _reservation_station_25_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_25_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_25_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_25_io_i_uop_valid = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_pc = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_inst = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_func_code = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_target = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_branch_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_select = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_taken = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_phy_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_stale_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_arch_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_inst_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_regWen = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_src1_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_phy_rs1 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_arch_rs1 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_src2_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_phy_rs2 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_arch_rs2 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_rob_idx = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_imm = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_src1_value = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_src2_value = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_op1_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_op2_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_alu_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_mem_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_25_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_25_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_25_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_25_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_26_clock = clock;
  assign reservation_station_26_reset = reset;
  assign reservation_station_26_io_i_issue_granted = (_issue1_func_code_T_26 | _io_o_issue_packs_1_T_26) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_26_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_26_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_26_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_26_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_26_io_i_write_slot = _reservation_station_26_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_26_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_26_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_26_io_i_uop_valid = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_pc = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_inst = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_func_code = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_target = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_branch_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_select = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_taken = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_phy_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_stale_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_arch_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_inst_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_regWen = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_src1_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_phy_rs1 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_arch_rs1 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_src2_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_phy_rs2 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_arch_rs2 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_rob_idx = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_imm = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_src1_value = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_src2_value = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_op1_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_op2_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_alu_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_mem_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_26_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_26_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_26_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_26_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_27_clock = clock;
  assign reservation_station_27_reset = reset;
  assign reservation_station_27_io_i_issue_granted = (_issue1_func_code_T_27 | _io_o_issue_packs_1_T_27) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_27_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_27_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_27_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_27_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_27_io_i_write_slot = _reservation_station_27_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_27_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_27_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_27_io_i_uop_valid = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_pc = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_inst = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_func_code = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_target = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_branch_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_select = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_taken = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_phy_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_stale_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_arch_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_inst_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_regWen = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_src1_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_phy_rs1 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_arch_rs1 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_src2_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_phy_rs2 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_arch_rs2 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_rob_idx = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_imm = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_src1_value = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_src2_value = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_op1_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_op2_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_alu_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_mem_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_27_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_27_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_27_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_27_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_28_clock = clock;
  assign reservation_station_28_reset = reset;
  assign reservation_station_28_io_i_issue_granted = (_issue1_func_code_T_28 | _io_o_issue_packs_1_T_28) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_28_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_28_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_28_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_28_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_28_io_i_write_slot = _reservation_station_28_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_28_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_28_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_28_io_i_uop_valid = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_pc = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_inst = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_func_code = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_target = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_branch_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_select = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_taken = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_phy_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_stale_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_arch_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_inst_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_regWen = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_src1_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_phy_rs1 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_arch_rs1 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_src2_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_phy_rs2 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_arch_rs2 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_rob_idx = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_imm = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_src1_value = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_src2_value = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_op1_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_op2_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_alu_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_mem_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_28_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_28_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_28_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_28_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_29_clock = clock;
  assign reservation_station_29_reset = reset;
  assign reservation_station_29_io_i_issue_granted = (_issue1_func_code_T_29 | _io_o_issue_packs_1_T_29) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_29_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_29_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_29_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_29_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_29_io_i_write_slot = _reservation_station_29_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_29_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_29_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_29_io_i_uop_valid = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_pc = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_inst = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_func_code = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_target = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_branch_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_select = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_taken = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_phy_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_stale_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_arch_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_inst_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_regWen = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_src1_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_phy_rs1 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_arch_rs1 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_src2_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_phy_rs2 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_arch_rs2 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_rob_idx = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_imm = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_src1_value = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_src2_value = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_op1_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_op2_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_alu_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_mem_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_29_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_29_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_29_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_29_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_30_clock = clock;
  assign reservation_station_30_reset = reset;
  assign reservation_station_30_io_i_issue_granted = (_issue1_func_code_T_30 | _io_o_issue_packs_1_T_30) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_30_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_30_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_30_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_30_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_30_io_i_write_slot = _reservation_station_30_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_30_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_30_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_30_io_i_uop_valid = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_pc = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_inst = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_func_code = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_target = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_branch_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_select = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_taken = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_phy_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_stale_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_arch_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_inst_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_regWen = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_src1_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_phy_rs1 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_arch_rs1 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_src2_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_phy_rs2 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_arch_rs2 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_rob_idx = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_imm = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_src1_value = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_src2_value = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_op1_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_op2_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_alu_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_mem_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_30_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_30_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_30_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_30_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_31_clock = clock;
  assign reservation_station_31_reset = reset;
  assign reservation_station_31_io_i_issue_granted = (_issue1_func_code_T_31 | _io_o_issue_packs_1_T_31) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_31_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_31_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_31_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_31_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_31_io_i_write_slot = _reservation_station_31_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_31_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_31_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_31_io_i_uop_valid = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_pc = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_inst = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_func_code = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_target = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_branch_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_select = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_taken = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_phy_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_stale_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_arch_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_inst_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_regWen = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_src1_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_phy_rs1 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_arch_rs1 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_src2_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_phy_rs2 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_arch_rs2 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_rob_idx = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_imm = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_src1_value = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_src2_value = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_op1_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_op2_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_alu_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_mem_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_31_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_31_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_31_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_31_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
endmodule

module Arch_RegFile(
  input  [63:0] io_i_pregs_0,
  input  [63:0] io_i_pregs_1,
  input  [63:0] io_i_pregs_2,
  input  [63:0] io_i_pregs_3,
  input  [63:0] io_i_pregs_4,
  input  [63:0] io_i_pregs_5,
  input  [63:0] io_i_pregs_6,
  input  [63:0] io_i_pregs_7,
  input  [63:0] io_i_pregs_8,
  input  [63:0] io_i_pregs_9,
  input  [63:0] io_i_pregs_10,
  input  [63:0] io_i_pregs_11,
  input  [63:0] io_i_pregs_12,
  input  [63:0] io_i_pregs_13,
  input  [63:0] io_i_pregs_14,
  input  [63:0] io_i_pregs_15,
  input  [63:0] io_i_pregs_16,
  input  [63:0] io_i_pregs_17,
  input  [63:0] io_i_pregs_18,
  input  [63:0] io_i_pregs_19,
  input  [63:0] io_i_pregs_20,
  input  [63:0] io_i_pregs_21,
  input  [63:0] io_i_pregs_22,
  input  [63:0] io_i_pregs_23,
  input  [63:0] io_i_pregs_24,
  input  [63:0] io_i_pregs_25,
  input  [63:0] io_i_pregs_26,
  input  [63:0] io_i_pregs_27,
  input  [63:0] io_i_pregs_28,
  input  [63:0] io_i_pregs_29,
  input  [63:0] io_i_pregs_30,
  input  [63:0] io_i_pregs_31,
  input  [63:0] io_i_pregs_32,
  input  [63:0] io_i_pregs_33,
  input  [63:0] io_i_pregs_34,
  input  [63:0] io_i_pregs_35,
  input  [63:0] io_i_pregs_36,
  input  [63:0] io_i_pregs_37,
  input  [63:0] io_i_pregs_38,
  input  [63:0] io_i_pregs_39,
  input  [63:0] io_i_pregs_40,
  input  [63:0] io_i_pregs_41,
  input  [63:0] io_i_pregs_42,
  input  [63:0] io_i_pregs_43,
  input  [63:0] io_i_pregs_44,
  input  [63:0] io_i_pregs_45,
  input  [63:0] io_i_pregs_46,
  input  [63:0] io_i_pregs_47,
  input  [63:0] io_i_pregs_48,
  input  [63:0] io_i_pregs_49,
  input  [63:0] io_i_pregs_50,
  input  [63:0] io_i_pregs_51,
  input  [63:0] io_i_pregs_52,
  input  [63:0] io_i_pregs_53,
  input  [63:0] io_i_pregs_54,
  input  [63:0] io_i_pregs_55,
  input  [63:0] io_i_pregs_56,
  input  [63:0] io_i_pregs_57,
  input  [63:0] io_i_pregs_58,
  input  [63:0] io_i_pregs_59,
  input  [63:0] io_i_pregs_60,
  input  [63:0] io_i_pregs_61,
  input  [63:0] io_i_pregs_62,
  input  [63:0] io_i_pregs_63,
  input  [63:0] io_i_pregs_64,
  input  [63:0] io_i_pregs_65,
  input  [63:0] io_i_pregs_66,
  input  [63:0] io_i_pregs_67,
  input  [63:0] io_i_pregs_68,
  input  [63:0] io_i_pregs_69,
  input  [63:0] io_i_pregs_70,
  input  [63:0] io_i_pregs_71,
  input  [63:0] io_i_pregs_72,
  input  [63:0] io_i_pregs_73,
  input  [63:0] io_i_pregs_74,
  input  [63:0] io_i_pregs_75,
  input  [63:0] io_i_pregs_76,
  input  [63:0] io_i_pregs_77,
  input  [63:0] io_i_pregs_78,
  input  [63:0] io_i_pregs_79,
  input  [63:0] io_i_pregs_80,
  input  [63:0] io_i_pregs_81,
  input  [63:0] io_i_pregs_82,
  input  [63:0] io_i_pregs_83,
  input  [63:0] io_i_pregs_84,
  input  [63:0] io_i_pregs_85,
  input  [63:0] io_i_pregs_86,
  input  [63:0] io_i_pregs_87,
  input  [63:0] io_i_pregs_88,
  input  [63:0] io_i_pregs_89,
  input  [63:0] io_i_pregs_90,
  input  [63:0] io_i_pregs_91,
  input  [63:0] io_i_pregs_92,
  input  [63:0] io_i_pregs_93,
  input  [63:0] io_i_pregs_94,
  input  [63:0] io_i_pregs_95,
  input  [63:0] io_i_pregs_96,
  input  [63:0] io_i_pregs_97,
  input  [63:0] io_i_pregs_98,
  input  [63:0] io_i_pregs_99,
  input  [63:0] io_i_pregs_100,
  input  [63:0] io_i_pregs_101,
  input  [63:0] io_i_pregs_102,
  input  [63:0] io_i_pregs_103,
  input  [63:0] io_i_pregs_104,
  input  [63:0] io_i_pregs_105,
  input  [63:0] io_i_pregs_106,
  input  [63:0] io_i_pregs_107,
  input  [63:0] io_i_pregs_108,
  input  [63:0] io_i_pregs_109,
  input  [63:0] io_i_pregs_110,
  input  [63:0] io_i_pregs_111,
  input  [63:0] io_i_pregs_112,
  input  [63:0] io_i_pregs_113,
  input  [63:0] io_i_pregs_114,
  input  [63:0] io_i_pregs_115,
  input  [63:0] io_i_pregs_116,
  input  [63:0] io_i_pregs_117,
  input  [63:0] io_i_pregs_118,
  input  [63:0] io_i_pregs_119,
  input  [63:0] io_i_pregs_120,
  input  [63:0] io_i_pregs_121,
  input  [63:0] io_i_pregs_122,
  input  [63:0] io_i_pregs_123,
  input  [63:0] io_i_pregs_124,
  input  [63:0] io_i_pregs_125,
  input  [63:0] io_i_pregs_126,
  input  [63:0] io_i_pregs_127,
  input  [6:0]  io_i_rename_table_0,
  input  [6:0]  io_i_rename_table_1,
  input  [6:0]  io_i_rename_table_2,
  input  [6:0]  io_i_rename_table_3,
  input  [6:0]  io_i_rename_table_4,
  input  [6:0]  io_i_rename_table_5,
  input  [6:0]  io_i_rename_table_6,
  input  [6:0]  io_i_rename_table_7,
  input  [6:0]  io_i_rename_table_8,
  input  [6:0]  io_i_rename_table_9,
  input  [6:0]  io_i_rename_table_10,
  input  [6:0]  io_i_rename_table_11,
  input  [6:0]  io_i_rename_table_12,
  input  [6:0]  io_i_rename_table_13,
  input  [6:0]  io_i_rename_table_14,
  input  [6:0]  io_i_rename_table_15,
  input  [6:0]  io_i_rename_table_16,
  input  [6:0]  io_i_rename_table_17,
  input  [6:0]  io_i_rename_table_18,
  input  [6:0]  io_i_rename_table_19,
  input  [6:0]  io_i_rename_table_20,
  input  [6:0]  io_i_rename_table_21,
  input  [6:0]  io_i_rename_table_22,
  input  [6:0]  io_i_rename_table_23,
  input  [6:0]  io_i_rename_table_24,
  input  [6:0]  io_i_rename_table_25,
  input  [6:0]  io_i_rename_table_26,
  input  [6:0]  io_i_rename_table_27,
  input  [6:0]  io_i_rename_table_28,
  input  [6:0]  io_i_rename_table_29,
  input  [6:0]  io_i_rename_table_30,
  input  [6:0]  io_i_rename_table_31,
  input  [63:0] io_i_csrs_0,
  input  [63:0] io_i_csrs_1,
  input  [63:0] io_i_csrs_2,
  input  [63:0] io_i_csrs_3,
  output [63:0] io_o_arch_regs_0,
  output [63:0] io_o_arch_regs_1,
  output [63:0] io_o_arch_regs_2,
  output [63:0] io_o_arch_regs_3,
  output [63:0] io_o_arch_regs_4,
  output [63:0] io_o_arch_regs_5,
  output [63:0] io_o_arch_regs_6,
  output [63:0] io_o_arch_regs_7,
  output [63:0] io_o_arch_regs_8,
  output [63:0] io_o_arch_regs_9,
  output [63:0] io_o_arch_regs_10,
  output [63:0] io_o_arch_regs_11,
  output [63:0] io_o_arch_regs_12,
  output [63:0] io_o_arch_regs_13,
  output [63:0] io_o_arch_regs_14,
  output [63:0] io_o_arch_regs_15,
  output [63:0] io_o_arch_regs_16,
  output [63:0] io_o_arch_regs_17,
  output [63:0] io_o_arch_regs_18,
  output [63:0] io_o_arch_regs_19,
  output [63:0] io_o_arch_regs_20,
  output [63:0] io_o_arch_regs_21,
  output [63:0] io_o_arch_regs_22,
  output [63:0] io_o_arch_regs_23,
  output [63:0] io_o_arch_regs_24,
  output [63:0] io_o_arch_regs_25,
  output [63:0] io_o_arch_regs_26,
  output [63:0] io_o_arch_regs_27,
  output [63:0] io_o_arch_regs_28,
  output [63:0] io_o_arch_regs_29,
  output [63:0] io_o_arch_regs_30,
  output [63:0] io_o_arch_regs_31,
  output [63:0] io_o_csr_regs_0,
  output [63:0] io_o_csr_regs_1,
  output [63:0] io_o_csr_regs_2,
  output [63:0] io_o_csr_regs_3
);
  wire [63:0] _GEN_1 = 7'h1 == io_i_rename_table_0 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2 = 7'h2 == io_i_rename_table_0 ? io_i_pregs_2 : _GEN_1; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3 = 7'h3 == io_i_rename_table_0 ? io_i_pregs_3 : _GEN_2; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4 = 7'h4 == io_i_rename_table_0 ? io_i_pregs_4 : _GEN_3; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_5 = 7'h5 == io_i_rename_table_0 ? io_i_pregs_5 : _GEN_4; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_6 = 7'h6 == io_i_rename_table_0 ? io_i_pregs_6 : _GEN_5; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_7 = 7'h7 == io_i_rename_table_0 ? io_i_pregs_7 : _GEN_6; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_8 = 7'h8 == io_i_rename_table_0 ? io_i_pregs_8 : _GEN_7; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_9 = 7'h9 == io_i_rename_table_0 ? io_i_pregs_9 : _GEN_8; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_10 = 7'ha == io_i_rename_table_0 ? io_i_pregs_10 : _GEN_9; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_11 = 7'hb == io_i_rename_table_0 ? io_i_pregs_11 : _GEN_10; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_12 = 7'hc == io_i_rename_table_0 ? io_i_pregs_12 : _GEN_11; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_13 = 7'hd == io_i_rename_table_0 ? io_i_pregs_13 : _GEN_12; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_14 = 7'he == io_i_rename_table_0 ? io_i_pregs_14 : _GEN_13; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_15 = 7'hf == io_i_rename_table_0 ? io_i_pregs_15 : _GEN_14; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_16 = 7'h10 == io_i_rename_table_0 ? io_i_pregs_16 : _GEN_15; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_17 = 7'h11 == io_i_rename_table_0 ? io_i_pregs_17 : _GEN_16; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_18 = 7'h12 == io_i_rename_table_0 ? io_i_pregs_18 : _GEN_17; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_19 = 7'h13 == io_i_rename_table_0 ? io_i_pregs_19 : _GEN_18; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_20 = 7'h14 == io_i_rename_table_0 ? io_i_pregs_20 : _GEN_19; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_21 = 7'h15 == io_i_rename_table_0 ? io_i_pregs_21 : _GEN_20; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_22 = 7'h16 == io_i_rename_table_0 ? io_i_pregs_22 : _GEN_21; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_23 = 7'h17 == io_i_rename_table_0 ? io_i_pregs_23 : _GEN_22; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_24 = 7'h18 == io_i_rename_table_0 ? io_i_pregs_24 : _GEN_23; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_25 = 7'h19 == io_i_rename_table_0 ? io_i_pregs_25 : _GEN_24; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_26 = 7'h1a == io_i_rename_table_0 ? io_i_pregs_26 : _GEN_25; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_27 = 7'h1b == io_i_rename_table_0 ? io_i_pregs_27 : _GEN_26; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_28 = 7'h1c == io_i_rename_table_0 ? io_i_pregs_28 : _GEN_27; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_29 = 7'h1d == io_i_rename_table_0 ? io_i_pregs_29 : _GEN_28; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_30 = 7'h1e == io_i_rename_table_0 ? io_i_pregs_30 : _GEN_29; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_31 = 7'h1f == io_i_rename_table_0 ? io_i_pregs_31 : _GEN_30; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_32 = 7'h20 == io_i_rename_table_0 ? io_i_pregs_32 : _GEN_31; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_33 = 7'h21 == io_i_rename_table_0 ? io_i_pregs_33 : _GEN_32; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_34 = 7'h22 == io_i_rename_table_0 ? io_i_pregs_34 : _GEN_33; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_35 = 7'h23 == io_i_rename_table_0 ? io_i_pregs_35 : _GEN_34; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_36 = 7'h24 == io_i_rename_table_0 ? io_i_pregs_36 : _GEN_35; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_37 = 7'h25 == io_i_rename_table_0 ? io_i_pregs_37 : _GEN_36; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_38 = 7'h26 == io_i_rename_table_0 ? io_i_pregs_38 : _GEN_37; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_39 = 7'h27 == io_i_rename_table_0 ? io_i_pregs_39 : _GEN_38; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_40 = 7'h28 == io_i_rename_table_0 ? io_i_pregs_40 : _GEN_39; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_41 = 7'h29 == io_i_rename_table_0 ? io_i_pregs_41 : _GEN_40; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_42 = 7'h2a == io_i_rename_table_0 ? io_i_pregs_42 : _GEN_41; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_43 = 7'h2b == io_i_rename_table_0 ? io_i_pregs_43 : _GEN_42; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_44 = 7'h2c == io_i_rename_table_0 ? io_i_pregs_44 : _GEN_43; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_45 = 7'h2d == io_i_rename_table_0 ? io_i_pregs_45 : _GEN_44; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_46 = 7'h2e == io_i_rename_table_0 ? io_i_pregs_46 : _GEN_45; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_47 = 7'h2f == io_i_rename_table_0 ? io_i_pregs_47 : _GEN_46; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_48 = 7'h30 == io_i_rename_table_0 ? io_i_pregs_48 : _GEN_47; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_49 = 7'h31 == io_i_rename_table_0 ? io_i_pregs_49 : _GEN_48; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_50 = 7'h32 == io_i_rename_table_0 ? io_i_pregs_50 : _GEN_49; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_51 = 7'h33 == io_i_rename_table_0 ? io_i_pregs_51 : _GEN_50; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_52 = 7'h34 == io_i_rename_table_0 ? io_i_pregs_52 : _GEN_51; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_53 = 7'h35 == io_i_rename_table_0 ? io_i_pregs_53 : _GEN_52; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_54 = 7'h36 == io_i_rename_table_0 ? io_i_pregs_54 : _GEN_53; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_55 = 7'h37 == io_i_rename_table_0 ? io_i_pregs_55 : _GEN_54; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_56 = 7'h38 == io_i_rename_table_0 ? io_i_pregs_56 : _GEN_55; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_57 = 7'h39 == io_i_rename_table_0 ? io_i_pregs_57 : _GEN_56; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_58 = 7'h3a == io_i_rename_table_0 ? io_i_pregs_58 : _GEN_57; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_59 = 7'h3b == io_i_rename_table_0 ? io_i_pregs_59 : _GEN_58; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_60 = 7'h3c == io_i_rename_table_0 ? io_i_pregs_60 : _GEN_59; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_61 = 7'h3d == io_i_rename_table_0 ? io_i_pregs_61 : _GEN_60; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_62 = 7'h3e == io_i_rename_table_0 ? io_i_pregs_62 : _GEN_61; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_63 = 7'h3f == io_i_rename_table_0 ? io_i_pregs_63 : _GEN_62; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_64 = 7'h40 == io_i_rename_table_0 ? io_i_pregs_64 : _GEN_63; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_65 = 7'h41 == io_i_rename_table_0 ? io_i_pregs_65 : _GEN_64; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_66 = 7'h42 == io_i_rename_table_0 ? io_i_pregs_66 : _GEN_65; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_67 = 7'h43 == io_i_rename_table_0 ? io_i_pregs_67 : _GEN_66; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_68 = 7'h44 == io_i_rename_table_0 ? io_i_pregs_68 : _GEN_67; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_69 = 7'h45 == io_i_rename_table_0 ? io_i_pregs_69 : _GEN_68; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_70 = 7'h46 == io_i_rename_table_0 ? io_i_pregs_70 : _GEN_69; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_71 = 7'h47 == io_i_rename_table_0 ? io_i_pregs_71 : _GEN_70; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_72 = 7'h48 == io_i_rename_table_0 ? io_i_pregs_72 : _GEN_71; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_73 = 7'h49 == io_i_rename_table_0 ? io_i_pregs_73 : _GEN_72; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_74 = 7'h4a == io_i_rename_table_0 ? io_i_pregs_74 : _GEN_73; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_75 = 7'h4b == io_i_rename_table_0 ? io_i_pregs_75 : _GEN_74; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_76 = 7'h4c == io_i_rename_table_0 ? io_i_pregs_76 : _GEN_75; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_77 = 7'h4d == io_i_rename_table_0 ? io_i_pregs_77 : _GEN_76; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_78 = 7'h4e == io_i_rename_table_0 ? io_i_pregs_78 : _GEN_77; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_79 = 7'h4f == io_i_rename_table_0 ? io_i_pregs_79 : _GEN_78; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_80 = 7'h50 == io_i_rename_table_0 ? io_i_pregs_80 : _GEN_79; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_81 = 7'h51 == io_i_rename_table_0 ? io_i_pregs_81 : _GEN_80; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_82 = 7'h52 == io_i_rename_table_0 ? io_i_pregs_82 : _GEN_81; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_83 = 7'h53 == io_i_rename_table_0 ? io_i_pregs_83 : _GEN_82; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_84 = 7'h54 == io_i_rename_table_0 ? io_i_pregs_84 : _GEN_83; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_85 = 7'h55 == io_i_rename_table_0 ? io_i_pregs_85 : _GEN_84; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_86 = 7'h56 == io_i_rename_table_0 ? io_i_pregs_86 : _GEN_85; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_87 = 7'h57 == io_i_rename_table_0 ? io_i_pregs_87 : _GEN_86; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_88 = 7'h58 == io_i_rename_table_0 ? io_i_pregs_88 : _GEN_87; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_89 = 7'h59 == io_i_rename_table_0 ? io_i_pregs_89 : _GEN_88; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_90 = 7'h5a == io_i_rename_table_0 ? io_i_pregs_90 : _GEN_89; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_91 = 7'h5b == io_i_rename_table_0 ? io_i_pregs_91 : _GEN_90; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_92 = 7'h5c == io_i_rename_table_0 ? io_i_pregs_92 : _GEN_91; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_93 = 7'h5d == io_i_rename_table_0 ? io_i_pregs_93 : _GEN_92; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_94 = 7'h5e == io_i_rename_table_0 ? io_i_pregs_94 : _GEN_93; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_95 = 7'h5f == io_i_rename_table_0 ? io_i_pregs_95 : _GEN_94; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_96 = 7'h60 == io_i_rename_table_0 ? io_i_pregs_96 : _GEN_95; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_97 = 7'h61 == io_i_rename_table_0 ? io_i_pregs_97 : _GEN_96; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_98 = 7'h62 == io_i_rename_table_0 ? io_i_pregs_98 : _GEN_97; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_99 = 7'h63 == io_i_rename_table_0 ? io_i_pregs_99 : _GEN_98; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_100 = 7'h64 == io_i_rename_table_0 ? io_i_pregs_100 : _GEN_99; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_101 = 7'h65 == io_i_rename_table_0 ? io_i_pregs_101 : _GEN_100; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_102 = 7'h66 == io_i_rename_table_0 ? io_i_pregs_102 : _GEN_101; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_103 = 7'h67 == io_i_rename_table_0 ? io_i_pregs_103 : _GEN_102; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_104 = 7'h68 == io_i_rename_table_0 ? io_i_pregs_104 : _GEN_103; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_105 = 7'h69 == io_i_rename_table_0 ? io_i_pregs_105 : _GEN_104; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_106 = 7'h6a == io_i_rename_table_0 ? io_i_pregs_106 : _GEN_105; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_107 = 7'h6b == io_i_rename_table_0 ? io_i_pregs_107 : _GEN_106; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_108 = 7'h6c == io_i_rename_table_0 ? io_i_pregs_108 : _GEN_107; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_109 = 7'h6d == io_i_rename_table_0 ? io_i_pregs_109 : _GEN_108; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_110 = 7'h6e == io_i_rename_table_0 ? io_i_pregs_110 : _GEN_109; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_111 = 7'h6f == io_i_rename_table_0 ? io_i_pregs_111 : _GEN_110; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_112 = 7'h70 == io_i_rename_table_0 ? io_i_pregs_112 : _GEN_111; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_113 = 7'h71 == io_i_rename_table_0 ? io_i_pregs_113 : _GEN_112; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_114 = 7'h72 == io_i_rename_table_0 ? io_i_pregs_114 : _GEN_113; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_115 = 7'h73 == io_i_rename_table_0 ? io_i_pregs_115 : _GEN_114; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_116 = 7'h74 == io_i_rename_table_0 ? io_i_pregs_116 : _GEN_115; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_117 = 7'h75 == io_i_rename_table_0 ? io_i_pregs_117 : _GEN_116; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_118 = 7'h76 == io_i_rename_table_0 ? io_i_pregs_118 : _GEN_117; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_119 = 7'h77 == io_i_rename_table_0 ? io_i_pregs_119 : _GEN_118; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_120 = 7'h78 == io_i_rename_table_0 ? io_i_pregs_120 : _GEN_119; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_121 = 7'h79 == io_i_rename_table_0 ? io_i_pregs_121 : _GEN_120; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_122 = 7'h7a == io_i_rename_table_0 ? io_i_pregs_122 : _GEN_121; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_123 = 7'h7b == io_i_rename_table_0 ? io_i_pregs_123 : _GEN_122; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_124 = 7'h7c == io_i_rename_table_0 ? io_i_pregs_124 : _GEN_123; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_125 = 7'h7d == io_i_rename_table_0 ? io_i_pregs_125 : _GEN_124; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_126 = 7'h7e == io_i_rename_table_0 ? io_i_pregs_126 : _GEN_125; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_129 = 7'h1 == io_i_rename_table_1 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_130 = 7'h2 == io_i_rename_table_1 ? io_i_pregs_2 : _GEN_129; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_131 = 7'h3 == io_i_rename_table_1 ? io_i_pregs_3 : _GEN_130; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_132 = 7'h4 == io_i_rename_table_1 ? io_i_pregs_4 : _GEN_131; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_133 = 7'h5 == io_i_rename_table_1 ? io_i_pregs_5 : _GEN_132; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_134 = 7'h6 == io_i_rename_table_1 ? io_i_pregs_6 : _GEN_133; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_135 = 7'h7 == io_i_rename_table_1 ? io_i_pregs_7 : _GEN_134; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_136 = 7'h8 == io_i_rename_table_1 ? io_i_pregs_8 : _GEN_135; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_137 = 7'h9 == io_i_rename_table_1 ? io_i_pregs_9 : _GEN_136; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_138 = 7'ha == io_i_rename_table_1 ? io_i_pregs_10 : _GEN_137; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_139 = 7'hb == io_i_rename_table_1 ? io_i_pregs_11 : _GEN_138; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_140 = 7'hc == io_i_rename_table_1 ? io_i_pregs_12 : _GEN_139; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_141 = 7'hd == io_i_rename_table_1 ? io_i_pregs_13 : _GEN_140; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_142 = 7'he == io_i_rename_table_1 ? io_i_pregs_14 : _GEN_141; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_143 = 7'hf == io_i_rename_table_1 ? io_i_pregs_15 : _GEN_142; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_144 = 7'h10 == io_i_rename_table_1 ? io_i_pregs_16 : _GEN_143; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_145 = 7'h11 == io_i_rename_table_1 ? io_i_pregs_17 : _GEN_144; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_146 = 7'h12 == io_i_rename_table_1 ? io_i_pregs_18 : _GEN_145; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_147 = 7'h13 == io_i_rename_table_1 ? io_i_pregs_19 : _GEN_146; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_148 = 7'h14 == io_i_rename_table_1 ? io_i_pregs_20 : _GEN_147; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_149 = 7'h15 == io_i_rename_table_1 ? io_i_pregs_21 : _GEN_148; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_150 = 7'h16 == io_i_rename_table_1 ? io_i_pregs_22 : _GEN_149; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_151 = 7'h17 == io_i_rename_table_1 ? io_i_pregs_23 : _GEN_150; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_152 = 7'h18 == io_i_rename_table_1 ? io_i_pregs_24 : _GEN_151; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_153 = 7'h19 == io_i_rename_table_1 ? io_i_pregs_25 : _GEN_152; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_154 = 7'h1a == io_i_rename_table_1 ? io_i_pregs_26 : _GEN_153; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_155 = 7'h1b == io_i_rename_table_1 ? io_i_pregs_27 : _GEN_154; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_156 = 7'h1c == io_i_rename_table_1 ? io_i_pregs_28 : _GEN_155; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_157 = 7'h1d == io_i_rename_table_1 ? io_i_pregs_29 : _GEN_156; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_158 = 7'h1e == io_i_rename_table_1 ? io_i_pregs_30 : _GEN_157; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_159 = 7'h1f == io_i_rename_table_1 ? io_i_pregs_31 : _GEN_158; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_160 = 7'h20 == io_i_rename_table_1 ? io_i_pregs_32 : _GEN_159; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_161 = 7'h21 == io_i_rename_table_1 ? io_i_pregs_33 : _GEN_160; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_162 = 7'h22 == io_i_rename_table_1 ? io_i_pregs_34 : _GEN_161; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_163 = 7'h23 == io_i_rename_table_1 ? io_i_pregs_35 : _GEN_162; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_164 = 7'h24 == io_i_rename_table_1 ? io_i_pregs_36 : _GEN_163; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_165 = 7'h25 == io_i_rename_table_1 ? io_i_pregs_37 : _GEN_164; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_166 = 7'h26 == io_i_rename_table_1 ? io_i_pregs_38 : _GEN_165; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_167 = 7'h27 == io_i_rename_table_1 ? io_i_pregs_39 : _GEN_166; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_168 = 7'h28 == io_i_rename_table_1 ? io_i_pregs_40 : _GEN_167; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_169 = 7'h29 == io_i_rename_table_1 ? io_i_pregs_41 : _GEN_168; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_170 = 7'h2a == io_i_rename_table_1 ? io_i_pregs_42 : _GEN_169; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_171 = 7'h2b == io_i_rename_table_1 ? io_i_pregs_43 : _GEN_170; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_172 = 7'h2c == io_i_rename_table_1 ? io_i_pregs_44 : _GEN_171; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_173 = 7'h2d == io_i_rename_table_1 ? io_i_pregs_45 : _GEN_172; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_174 = 7'h2e == io_i_rename_table_1 ? io_i_pregs_46 : _GEN_173; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_175 = 7'h2f == io_i_rename_table_1 ? io_i_pregs_47 : _GEN_174; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_176 = 7'h30 == io_i_rename_table_1 ? io_i_pregs_48 : _GEN_175; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_177 = 7'h31 == io_i_rename_table_1 ? io_i_pregs_49 : _GEN_176; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_178 = 7'h32 == io_i_rename_table_1 ? io_i_pregs_50 : _GEN_177; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_179 = 7'h33 == io_i_rename_table_1 ? io_i_pregs_51 : _GEN_178; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_180 = 7'h34 == io_i_rename_table_1 ? io_i_pregs_52 : _GEN_179; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_181 = 7'h35 == io_i_rename_table_1 ? io_i_pregs_53 : _GEN_180; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_182 = 7'h36 == io_i_rename_table_1 ? io_i_pregs_54 : _GEN_181; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_183 = 7'h37 == io_i_rename_table_1 ? io_i_pregs_55 : _GEN_182; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_184 = 7'h38 == io_i_rename_table_1 ? io_i_pregs_56 : _GEN_183; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_185 = 7'h39 == io_i_rename_table_1 ? io_i_pregs_57 : _GEN_184; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_186 = 7'h3a == io_i_rename_table_1 ? io_i_pregs_58 : _GEN_185; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_187 = 7'h3b == io_i_rename_table_1 ? io_i_pregs_59 : _GEN_186; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_188 = 7'h3c == io_i_rename_table_1 ? io_i_pregs_60 : _GEN_187; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_189 = 7'h3d == io_i_rename_table_1 ? io_i_pregs_61 : _GEN_188; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_190 = 7'h3e == io_i_rename_table_1 ? io_i_pregs_62 : _GEN_189; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_191 = 7'h3f == io_i_rename_table_1 ? io_i_pregs_63 : _GEN_190; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_192 = 7'h40 == io_i_rename_table_1 ? io_i_pregs_64 : _GEN_191; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_193 = 7'h41 == io_i_rename_table_1 ? io_i_pregs_65 : _GEN_192; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_194 = 7'h42 == io_i_rename_table_1 ? io_i_pregs_66 : _GEN_193; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_195 = 7'h43 == io_i_rename_table_1 ? io_i_pregs_67 : _GEN_194; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_196 = 7'h44 == io_i_rename_table_1 ? io_i_pregs_68 : _GEN_195; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_197 = 7'h45 == io_i_rename_table_1 ? io_i_pregs_69 : _GEN_196; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_198 = 7'h46 == io_i_rename_table_1 ? io_i_pregs_70 : _GEN_197; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_199 = 7'h47 == io_i_rename_table_1 ? io_i_pregs_71 : _GEN_198; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_200 = 7'h48 == io_i_rename_table_1 ? io_i_pregs_72 : _GEN_199; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_201 = 7'h49 == io_i_rename_table_1 ? io_i_pregs_73 : _GEN_200; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_202 = 7'h4a == io_i_rename_table_1 ? io_i_pregs_74 : _GEN_201; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_203 = 7'h4b == io_i_rename_table_1 ? io_i_pregs_75 : _GEN_202; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_204 = 7'h4c == io_i_rename_table_1 ? io_i_pregs_76 : _GEN_203; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_205 = 7'h4d == io_i_rename_table_1 ? io_i_pregs_77 : _GEN_204; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_206 = 7'h4e == io_i_rename_table_1 ? io_i_pregs_78 : _GEN_205; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_207 = 7'h4f == io_i_rename_table_1 ? io_i_pregs_79 : _GEN_206; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_208 = 7'h50 == io_i_rename_table_1 ? io_i_pregs_80 : _GEN_207; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_209 = 7'h51 == io_i_rename_table_1 ? io_i_pregs_81 : _GEN_208; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_210 = 7'h52 == io_i_rename_table_1 ? io_i_pregs_82 : _GEN_209; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_211 = 7'h53 == io_i_rename_table_1 ? io_i_pregs_83 : _GEN_210; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_212 = 7'h54 == io_i_rename_table_1 ? io_i_pregs_84 : _GEN_211; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_213 = 7'h55 == io_i_rename_table_1 ? io_i_pregs_85 : _GEN_212; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_214 = 7'h56 == io_i_rename_table_1 ? io_i_pregs_86 : _GEN_213; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_215 = 7'h57 == io_i_rename_table_1 ? io_i_pregs_87 : _GEN_214; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_216 = 7'h58 == io_i_rename_table_1 ? io_i_pregs_88 : _GEN_215; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_217 = 7'h59 == io_i_rename_table_1 ? io_i_pregs_89 : _GEN_216; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_218 = 7'h5a == io_i_rename_table_1 ? io_i_pregs_90 : _GEN_217; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_219 = 7'h5b == io_i_rename_table_1 ? io_i_pregs_91 : _GEN_218; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_220 = 7'h5c == io_i_rename_table_1 ? io_i_pregs_92 : _GEN_219; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_221 = 7'h5d == io_i_rename_table_1 ? io_i_pregs_93 : _GEN_220; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_222 = 7'h5e == io_i_rename_table_1 ? io_i_pregs_94 : _GEN_221; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_223 = 7'h5f == io_i_rename_table_1 ? io_i_pregs_95 : _GEN_222; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_224 = 7'h60 == io_i_rename_table_1 ? io_i_pregs_96 : _GEN_223; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_225 = 7'h61 == io_i_rename_table_1 ? io_i_pregs_97 : _GEN_224; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_226 = 7'h62 == io_i_rename_table_1 ? io_i_pregs_98 : _GEN_225; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_227 = 7'h63 == io_i_rename_table_1 ? io_i_pregs_99 : _GEN_226; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_228 = 7'h64 == io_i_rename_table_1 ? io_i_pregs_100 : _GEN_227; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_229 = 7'h65 == io_i_rename_table_1 ? io_i_pregs_101 : _GEN_228; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_230 = 7'h66 == io_i_rename_table_1 ? io_i_pregs_102 : _GEN_229; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_231 = 7'h67 == io_i_rename_table_1 ? io_i_pregs_103 : _GEN_230; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_232 = 7'h68 == io_i_rename_table_1 ? io_i_pregs_104 : _GEN_231; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_233 = 7'h69 == io_i_rename_table_1 ? io_i_pregs_105 : _GEN_232; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_234 = 7'h6a == io_i_rename_table_1 ? io_i_pregs_106 : _GEN_233; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_235 = 7'h6b == io_i_rename_table_1 ? io_i_pregs_107 : _GEN_234; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_236 = 7'h6c == io_i_rename_table_1 ? io_i_pregs_108 : _GEN_235; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_237 = 7'h6d == io_i_rename_table_1 ? io_i_pregs_109 : _GEN_236; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_238 = 7'h6e == io_i_rename_table_1 ? io_i_pregs_110 : _GEN_237; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_239 = 7'h6f == io_i_rename_table_1 ? io_i_pregs_111 : _GEN_238; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_240 = 7'h70 == io_i_rename_table_1 ? io_i_pregs_112 : _GEN_239; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_241 = 7'h71 == io_i_rename_table_1 ? io_i_pregs_113 : _GEN_240; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_242 = 7'h72 == io_i_rename_table_1 ? io_i_pregs_114 : _GEN_241; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_243 = 7'h73 == io_i_rename_table_1 ? io_i_pregs_115 : _GEN_242; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_244 = 7'h74 == io_i_rename_table_1 ? io_i_pregs_116 : _GEN_243; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_245 = 7'h75 == io_i_rename_table_1 ? io_i_pregs_117 : _GEN_244; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_246 = 7'h76 == io_i_rename_table_1 ? io_i_pregs_118 : _GEN_245; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_247 = 7'h77 == io_i_rename_table_1 ? io_i_pregs_119 : _GEN_246; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_248 = 7'h78 == io_i_rename_table_1 ? io_i_pregs_120 : _GEN_247; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_249 = 7'h79 == io_i_rename_table_1 ? io_i_pregs_121 : _GEN_248; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_250 = 7'h7a == io_i_rename_table_1 ? io_i_pregs_122 : _GEN_249; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_251 = 7'h7b == io_i_rename_table_1 ? io_i_pregs_123 : _GEN_250; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_252 = 7'h7c == io_i_rename_table_1 ? io_i_pregs_124 : _GEN_251; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_253 = 7'h7d == io_i_rename_table_1 ? io_i_pregs_125 : _GEN_252; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_254 = 7'h7e == io_i_rename_table_1 ? io_i_pregs_126 : _GEN_253; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_257 = 7'h1 == io_i_rename_table_2 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_258 = 7'h2 == io_i_rename_table_2 ? io_i_pregs_2 : _GEN_257; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_259 = 7'h3 == io_i_rename_table_2 ? io_i_pregs_3 : _GEN_258; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_260 = 7'h4 == io_i_rename_table_2 ? io_i_pregs_4 : _GEN_259; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_261 = 7'h5 == io_i_rename_table_2 ? io_i_pregs_5 : _GEN_260; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_262 = 7'h6 == io_i_rename_table_2 ? io_i_pregs_6 : _GEN_261; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_263 = 7'h7 == io_i_rename_table_2 ? io_i_pregs_7 : _GEN_262; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_264 = 7'h8 == io_i_rename_table_2 ? io_i_pregs_8 : _GEN_263; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_265 = 7'h9 == io_i_rename_table_2 ? io_i_pregs_9 : _GEN_264; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_266 = 7'ha == io_i_rename_table_2 ? io_i_pregs_10 : _GEN_265; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_267 = 7'hb == io_i_rename_table_2 ? io_i_pregs_11 : _GEN_266; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_268 = 7'hc == io_i_rename_table_2 ? io_i_pregs_12 : _GEN_267; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_269 = 7'hd == io_i_rename_table_2 ? io_i_pregs_13 : _GEN_268; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_270 = 7'he == io_i_rename_table_2 ? io_i_pregs_14 : _GEN_269; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_271 = 7'hf == io_i_rename_table_2 ? io_i_pregs_15 : _GEN_270; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_272 = 7'h10 == io_i_rename_table_2 ? io_i_pregs_16 : _GEN_271; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_273 = 7'h11 == io_i_rename_table_2 ? io_i_pregs_17 : _GEN_272; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_274 = 7'h12 == io_i_rename_table_2 ? io_i_pregs_18 : _GEN_273; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_275 = 7'h13 == io_i_rename_table_2 ? io_i_pregs_19 : _GEN_274; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_276 = 7'h14 == io_i_rename_table_2 ? io_i_pregs_20 : _GEN_275; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_277 = 7'h15 == io_i_rename_table_2 ? io_i_pregs_21 : _GEN_276; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_278 = 7'h16 == io_i_rename_table_2 ? io_i_pregs_22 : _GEN_277; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_279 = 7'h17 == io_i_rename_table_2 ? io_i_pregs_23 : _GEN_278; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_280 = 7'h18 == io_i_rename_table_2 ? io_i_pregs_24 : _GEN_279; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_281 = 7'h19 == io_i_rename_table_2 ? io_i_pregs_25 : _GEN_280; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_282 = 7'h1a == io_i_rename_table_2 ? io_i_pregs_26 : _GEN_281; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_283 = 7'h1b == io_i_rename_table_2 ? io_i_pregs_27 : _GEN_282; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_284 = 7'h1c == io_i_rename_table_2 ? io_i_pregs_28 : _GEN_283; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_285 = 7'h1d == io_i_rename_table_2 ? io_i_pregs_29 : _GEN_284; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_286 = 7'h1e == io_i_rename_table_2 ? io_i_pregs_30 : _GEN_285; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_287 = 7'h1f == io_i_rename_table_2 ? io_i_pregs_31 : _GEN_286; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_288 = 7'h20 == io_i_rename_table_2 ? io_i_pregs_32 : _GEN_287; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_289 = 7'h21 == io_i_rename_table_2 ? io_i_pregs_33 : _GEN_288; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_290 = 7'h22 == io_i_rename_table_2 ? io_i_pregs_34 : _GEN_289; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_291 = 7'h23 == io_i_rename_table_2 ? io_i_pregs_35 : _GEN_290; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_292 = 7'h24 == io_i_rename_table_2 ? io_i_pregs_36 : _GEN_291; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_293 = 7'h25 == io_i_rename_table_2 ? io_i_pregs_37 : _GEN_292; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_294 = 7'h26 == io_i_rename_table_2 ? io_i_pregs_38 : _GEN_293; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_295 = 7'h27 == io_i_rename_table_2 ? io_i_pregs_39 : _GEN_294; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_296 = 7'h28 == io_i_rename_table_2 ? io_i_pregs_40 : _GEN_295; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_297 = 7'h29 == io_i_rename_table_2 ? io_i_pregs_41 : _GEN_296; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_298 = 7'h2a == io_i_rename_table_2 ? io_i_pregs_42 : _GEN_297; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_299 = 7'h2b == io_i_rename_table_2 ? io_i_pregs_43 : _GEN_298; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_300 = 7'h2c == io_i_rename_table_2 ? io_i_pregs_44 : _GEN_299; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_301 = 7'h2d == io_i_rename_table_2 ? io_i_pregs_45 : _GEN_300; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_302 = 7'h2e == io_i_rename_table_2 ? io_i_pregs_46 : _GEN_301; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_303 = 7'h2f == io_i_rename_table_2 ? io_i_pregs_47 : _GEN_302; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_304 = 7'h30 == io_i_rename_table_2 ? io_i_pregs_48 : _GEN_303; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_305 = 7'h31 == io_i_rename_table_2 ? io_i_pregs_49 : _GEN_304; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_306 = 7'h32 == io_i_rename_table_2 ? io_i_pregs_50 : _GEN_305; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_307 = 7'h33 == io_i_rename_table_2 ? io_i_pregs_51 : _GEN_306; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_308 = 7'h34 == io_i_rename_table_2 ? io_i_pregs_52 : _GEN_307; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_309 = 7'h35 == io_i_rename_table_2 ? io_i_pregs_53 : _GEN_308; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_310 = 7'h36 == io_i_rename_table_2 ? io_i_pregs_54 : _GEN_309; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_311 = 7'h37 == io_i_rename_table_2 ? io_i_pregs_55 : _GEN_310; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_312 = 7'h38 == io_i_rename_table_2 ? io_i_pregs_56 : _GEN_311; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_313 = 7'h39 == io_i_rename_table_2 ? io_i_pregs_57 : _GEN_312; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_314 = 7'h3a == io_i_rename_table_2 ? io_i_pregs_58 : _GEN_313; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_315 = 7'h3b == io_i_rename_table_2 ? io_i_pregs_59 : _GEN_314; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_316 = 7'h3c == io_i_rename_table_2 ? io_i_pregs_60 : _GEN_315; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_317 = 7'h3d == io_i_rename_table_2 ? io_i_pregs_61 : _GEN_316; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_318 = 7'h3e == io_i_rename_table_2 ? io_i_pregs_62 : _GEN_317; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_319 = 7'h3f == io_i_rename_table_2 ? io_i_pregs_63 : _GEN_318; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_320 = 7'h40 == io_i_rename_table_2 ? io_i_pregs_64 : _GEN_319; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_321 = 7'h41 == io_i_rename_table_2 ? io_i_pregs_65 : _GEN_320; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_322 = 7'h42 == io_i_rename_table_2 ? io_i_pregs_66 : _GEN_321; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_323 = 7'h43 == io_i_rename_table_2 ? io_i_pregs_67 : _GEN_322; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_324 = 7'h44 == io_i_rename_table_2 ? io_i_pregs_68 : _GEN_323; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_325 = 7'h45 == io_i_rename_table_2 ? io_i_pregs_69 : _GEN_324; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_326 = 7'h46 == io_i_rename_table_2 ? io_i_pregs_70 : _GEN_325; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_327 = 7'h47 == io_i_rename_table_2 ? io_i_pregs_71 : _GEN_326; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_328 = 7'h48 == io_i_rename_table_2 ? io_i_pregs_72 : _GEN_327; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_329 = 7'h49 == io_i_rename_table_2 ? io_i_pregs_73 : _GEN_328; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_330 = 7'h4a == io_i_rename_table_2 ? io_i_pregs_74 : _GEN_329; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_331 = 7'h4b == io_i_rename_table_2 ? io_i_pregs_75 : _GEN_330; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_332 = 7'h4c == io_i_rename_table_2 ? io_i_pregs_76 : _GEN_331; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_333 = 7'h4d == io_i_rename_table_2 ? io_i_pregs_77 : _GEN_332; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_334 = 7'h4e == io_i_rename_table_2 ? io_i_pregs_78 : _GEN_333; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_335 = 7'h4f == io_i_rename_table_2 ? io_i_pregs_79 : _GEN_334; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_336 = 7'h50 == io_i_rename_table_2 ? io_i_pregs_80 : _GEN_335; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_337 = 7'h51 == io_i_rename_table_2 ? io_i_pregs_81 : _GEN_336; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_338 = 7'h52 == io_i_rename_table_2 ? io_i_pregs_82 : _GEN_337; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_339 = 7'h53 == io_i_rename_table_2 ? io_i_pregs_83 : _GEN_338; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_340 = 7'h54 == io_i_rename_table_2 ? io_i_pregs_84 : _GEN_339; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_341 = 7'h55 == io_i_rename_table_2 ? io_i_pregs_85 : _GEN_340; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_342 = 7'h56 == io_i_rename_table_2 ? io_i_pregs_86 : _GEN_341; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_343 = 7'h57 == io_i_rename_table_2 ? io_i_pregs_87 : _GEN_342; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_344 = 7'h58 == io_i_rename_table_2 ? io_i_pregs_88 : _GEN_343; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_345 = 7'h59 == io_i_rename_table_2 ? io_i_pregs_89 : _GEN_344; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_346 = 7'h5a == io_i_rename_table_2 ? io_i_pregs_90 : _GEN_345; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_347 = 7'h5b == io_i_rename_table_2 ? io_i_pregs_91 : _GEN_346; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_348 = 7'h5c == io_i_rename_table_2 ? io_i_pregs_92 : _GEN_347; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_349 = 7'h5d == io_i_rename_table_2 ? io_i_pregs_93 : _GEN_348; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_350 = 7'h5e == io_i_rename_table_2 ? io_i_pregs_94 : _GEN_349; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_351 = 7'h5f == io_i_rename_table_2 ? io_i_pregs_95 : _GEN_350; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_352 = 7'h60 == io_i_rename_table_2 ? io_i_pregs_96 : _GEN_351; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_353 = 7'h61 == io_i_rename_table_2 ? io_i_pregs_97 : _GEN_352; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_354 = 7'h62 == io_i_rename_table_2 ? io_i_pregs_98 : _GEN_353; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_355 = 7'h63 == io_i_rename_table_2 ? io_i_pregs_99 : _GEN_354; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_356 = 7'h64 == io_i_rename_table_2 ? io_i_pregs_100 : _GEN_355; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_357 = 7'h65 == io_i_rename_table_2 ? io_i_pregs_101 : _GEN_356; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_358 = 7'h66 == io_i_rename_table_2 ? io_i_pregs_102 : _GEN_357; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_359 = 7'h67 == io_i_rename_table_2 ? io_i_pregs_103 : _GEN_358; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_360 = 7'h68 == io_i_rename_table_2 ? io_i_pregs_104 : _GEN_359; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_361 = 7'h69 == io_i_rename_table_2 ? io_i_pregs_105 : _GEN_360; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_362 = 7'h6a == io_i_rename_table_2 ? io_i_pregs_106 : _GEN_361; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_363 = 7'h6b == io_i_rename_table_2 ? io_i_pregs_107 : _GEN_362; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_364 = 7'h6c == io_i_rename_table_2 ? io_i_pregs_108 : _GEN_363; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_365 = 7'h6d == io_i_rename_table_2 ? io_i_pregs_109 : _GEN_364; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_366 = 7'h6e == io_i_rename_table_2 ? io_i_pregs_110 : _GEN_365; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_367 = 7'h6f == io_i_rename_table_2 ? io_i_pregs_111 : _GEN_366; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_368 = 7'h70 == io_i_rename_table_2 ? io_i_pregs_112 : _GEN_367; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_369 = 7'h71 == io_i_rename_table_2 ? io_i_pregs_113 : _GEN_368; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_370 = 7'h72 == io_i_rename_table_2 ? io_i_pregs_114 : _GEN_369; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_371 = 7'h73 == io_i_rename_table_2 ? io_i_pregs_115 : _GEN_370; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_372 = 7'h74 == io_i_rename_table_2 ? io_i_pregs_116 : _GEN_371; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_373 = 7'h75 == io_i_rename_table_2 ? io_i_pregs_117 : _GEN_372; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_374 = 7'h76 == io_i_rename_table_2 ? io_i_pregs_118 : _GEN_373; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_375 = 7'h77 == io_i_rename_table_2 ? io_i_pregs_119 : _GEN_374; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_376 = 7'h78 == io_i_rename_table_2 ? io_i_pregs_120 : _GEN_375; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_377 = 7'h79 == io_i_rename_table_2 ? io_i_pregs_121 : _GEN_376; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_378 = 7'h7a == io_i_rename_table_2 ? io_i_pregs_122 : _GEN_377; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_379 = 7'h7b == io_i_rename_table_2 ? io_i_pregs_123 : _GEN_378; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_380 = 7'h7c == io_i_rename_table_2 ? io_i_pregs_124 : _GEN_379; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_381 = 7'h7d == io_i_rename_table_2 ? io_i_pregs_125 : _GEN_380; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_382 = 7'h7e == io_i_rename_table_2 ? io_i_pregs_126 : _GEN_381; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_385 = 7'h1 == io_i_rename_table_3 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_386 = 7'h2 == io_i_rename_table_3 ? io_i_pregs_2 : _GEN_385; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_387 = 7'h3 == io_i_rename_table_3 ? io_i_pregs_3 : _GEN_386; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_388 = 7'h4 == io_i_rename_table_3 ? io_i_pregs_4 : _GEN_387; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_389 = 7'h5 == io_i_rename_table_3 ? io_i_pregs_5 : _GEN_388; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_390 = 7'h6 == io_i_rename_table_3 ? io_i_pregs_6 : _GEN_389; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_391 = 7'h7 == io_i_rename_table_3 ? io_i_pregs_7 : _GEN_390; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_392 = 7'h8 == io_i_rename_table_3 ? io_i_pregs_8 : _GEN_391; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_393 = 7'h9 == io_i_rename_table_3 ? io_i_pregs_9 : _GEN_392; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_394 = 7'ha == io_i_rename_table_3 ? io_i_pregs_10 : _GEN_393; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_395 = 7'hb == io_i_rename_table_3 ? io_i_pregs_11 : _GEN_394; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_396 = 7'hc == io_i_rename_table_3 ? io_i_pregs_12 : _GEN_395; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_397 = 7'hd == io_i_rename_table_3 ? io_i_pregs_13 : _GEN_396; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_398 = 7'he == io_i_rename_table_3 ? io_i_pregs_14 : _GEN_397; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_399 = 7'hf == io_i_rename_table_3 ? io_i_pregs_15 : _GEN_398; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_400 = 7'h10 == io_i_rename_table_3 ? io_i_pregs_16 : _GEN_399; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_401 = 7'h11 == io_i_rename_table_3 ? io_i_pregs_17 : _GEN_400; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_402 = 7'h12 == io_i_rename_table_3 ? io_i_pregs_18 : _GEN_401; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_403 = 7'h13 == io_i_rename_table_3 ? io_i_pregs_19 : _GEN_402; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_404 = 7'h14 == io_i_rename_table_3 ? io_i_pregs_20 : _GEN_403; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_405 = 7'h15 == io_i_rename_table_3 ? io_i_pregs_21 : _GEN_404; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_406 = 7'h16 == io_i_rename_table_3 ? io_i_pregs_22 : _GEN_405; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_407 = 7'h17 == io_i_rename_table_3 ? io_i_pregs_23 : _GEN_406; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_408 = 7'h18 == io_i_rename_table_3 ? io_i_pregs_24 : _GEN_407; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_409 = 7'h19 == io_i_rename_table_3 ? io_i_pregs_25 : _GEN_408; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_410 = 7'h1a == io_i_rename_table_3 ? io_i_pregs_26 : _GEN_409; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_411 = 7'h1b == io_i_rename_table_3 ? io_i_pregs_27 : _GEN_410; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_412 = 7'h1c == io_i_rename_table_3 ? io_i_pregs_28 : _GEN_411; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_413 = 7'h1d == io_i_rename_table_3 ? io_i_pregs_29 : _GEN_412; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_414 = 7'h1e == io_i_rename_table_3 ? io_i_pregs_30 : _GEN_413; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_415 = 7'h1f == io_i_rename_table_3 ? io_i_pregs_31 : _GEN_414; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_416 = 7'h20 == io_i_rename_table_3 ? io_i_pregs_32 : _GEN_415; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_417 = 7'h21 == io_i_rename_table_3 ? io_i_pregs_33 : _GEN_416; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_418 = 7'h22 == io_i_rename_table_3 ? io_i_pregs_34 : _GEN_417; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_419 = 7'h23 == io_i_rename_table_3 ? io_i_pregs_35 : _GEN_418; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_420 = 7'h24 == io_i_rename_table_3 ? io_i_pregs_36 : _GEN_419; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_421 = 7'h25 == io_i_rename_table_3 ? io_i_pregs_37 : _GEN_420; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_422 = 7'h26 == io_i_rename_table_3 ? io_i_pregs_38 : _GEN_421; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_423 = 7'h27 == io_i_rename_table_3 ? io_i_pregs_39 : _GEN_422; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_424 = 7'h28 == io_i_rename_table_3 ? io_i_pregs_40 : _GEN_423; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_425 = 7'h29 == io_i_rename_table_3 ? io_i_pregs_41 : _GEN_424; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_426 = 7'h2a == io_i_rename_table_3 ? io_i_pregs_42 : _GEN_425; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_427 = 7'h2b == io_i_rename_table_3 ? io_i_pregs_43 : _GEN_426; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_428 = 7'h2c == io_i_rename_table_3 ? io_i_pregs_44 : _GEN_427; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_429 = 7'h2d == io_i_rename_table_3 ? io_i_pregs_45 : _GEN_428; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_430 = 7'h2e == io_i_rename_table_3 ? io_i_pregs_46 : _GEN_429; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_431 = 7'h2f == io_i_rename_table_3 ? io_i_pregs_47 : _GEN_430; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_432 = 7'h30 == io_i_rename_table_3 ? io_i_pregs_48 : _GEN_431; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_433 = 7'h31 == io_i_rename_table_3 ? io_i_pregs_49 : _GEN_432; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_434 = 7'h32 == io_i_rename_table_3 ? io_i_pregs_50 : _GEN_433; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_435 = 7'h33 == io_i_rename_table_3 ? io_i_pregs_51 : _GEN_434; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_436 = 7'h34 == io_i_rename_table_3 ? io_i_pregs_52 : _GEN_435; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_437 = 7'h35 == io_i_rename_table_3 ? io_i_pregs_53 : _GEN_436; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_438 = 7'h36 == io_i_rename_table_3 ? io_i_pregs_54 : _GEN_437; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_439 = 7'h37 == io_i_rename_table_3 ? io_i_pregs_55 : _GEN_438; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_440 = 7'h38 == io_i_rename_table_3 ? io_i_pregs_56 : _GEN_439; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_441 = 7'h39 == io_i_rename_table_3 ? io_i_pregs_57 : _GEN_440; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_442 = 7'h3a == io_i_rename_table_3 ? io_i_pregs_58 : _GEN_441; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_443 = 7'h3b == io_i_rename_table_3 ? io_i_pregs_59 : _GEN_442; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_444 = 7'h3c == io_i_rename_table_3 ? io_i_pregs_60 : _GEN_443; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_445 = 7'h3d == io_i_rename_table_3 ? io_i_pregs_61 : _GEN_444; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_446 = 7'h3e == io_i_rename_table_3 ? io_i_pregs_62 : _GEN_445; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_447 = 7'h3f == io_i_rename_table_3 ? io_i_pregs_63 : _GEN_446; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_448 = 7'h40 == io_i_rename_table_3 ? io_i_pregs_64 : _GEN_447; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_449 = 7'h41 == io_i_rename_table_3 ? io_i_pregs_65 : _GEN_448; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_450 = 7'h42 == io_i_rename_table_3 ? io_i_pregs_66 : _GEN_449; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_451 = 7'h43 == io_i_rename_table_3 ? io_i_pregs_67 : _GEN_450; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_452 = 7'h44 == io_i_rename_table_3 ? io_i_pregs_68 : _GEN_451; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_453 = 7'h45 == io_i_rename_table_3 ? io_i_pregs_69 : _GEN_452; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_454 = 7'h46 == io_i_rename_table_3 ? io_i_pregs_70 : _GEN_453; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_455 = 7'h47 == io_i_rename_table_3 ? io_i_pregs_71 : _GEN_454; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_456 = 7'h48 == io_i_rename_table_3 ? io_i_pregs_72 : _GEN_455; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_457 = 7'h49 == io_i_rename_table_3 ? io_i_pregs_73 : _GEN_456; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_458 = 7'h4a == io_i_rename_table_3 ? io_i_pregs_74 : _GEN_457; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_459 = 7'h4b == io_i_rename_table_3 ? io_i_pregs_75 : _GEN_458; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_460 = 7'h4c == io_i_rename_table_3 ? io_i_pregs_76 : _GEN_459; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_461 = 7'h4d == io_i_rename_table_3 ? io_i_pregs_77 : _GEN_460; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_462 = 7'h4e == io_i_rename_table_3 ? io_i_pregs_78 : _GEN_461; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_463 = 7'h4f == io_i_rename_table_3 ? io_i_pregs_79 : _GEN_462; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_464 = 7'h50 == io_i_rename_table_3 ? io_i_pregs_80 : _GEN_463; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_465 = 7'h51 == io_i_rename_table_3 ? io_i_pregs_81 : _GEN_464; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_466 = 7'h52 == io_i_rename_table_3 ? io_i_pregs_82 : _GEN_465; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_467 = 7'h53 == io_i_rename_table_3 ? io_i_pregs_83 : _GEN_466; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_468 = 7'h54 == io_i_rename_table_3 ? io_i_pregs_84 : _GEN_467; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_469 = 7'h55 == io_i_rename_table_3 ? io_i_pregs_85 : _GEN_468; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_470 = 7'h56 == io_i_rename_table_3 ? io_i_pregs_86 : _GEN_469; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_471 = 7'h57 == io_i_rename_table_3 ? io_i_pregs_87 : _GEN_470; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_472 = 7'h58 == io_i_rename_table_3 ? io_i_pregs_88 : _GEN_471; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_473 = 7'h59 == io_i_rename_table_3 ? io_i_pregs_89 : _GEN_472; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_474 = 7'h5a == io_i_rename_table_3 ? io_i_pregs_90 : _GEN_473; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_475 = 7'h5b == io_i_rename_table_3 ? io_i_pregs_91 : _GEN_474; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_476 = 7'h5c == io_i_rename_table_3 ? io_i_pregs_92 : _GEN_475; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_477 = 7'h5d == io_i_rename_table_3 ? io_i_pregs_93 : _GEN_476; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_478 = 7'h5e == io_i_rename_table_3 ? io_i_pregs_94 : _GEN_477; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_479 = 7'h5f == io_i_rename_table_3 ? io_i_pregs_95 : _GEN_478; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_480 = 7'h60 == io_i_rename_table_3 ? io_i_pregs_96 : _GEN_479; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_481 = 7'h61 == io_i_rename_table_3 ? io_i_pregs_97 : _GEN_480; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_482 = 7'h62 == io_i_rename_table_3 ? io_i_pregs_98 : _GEN_481; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_483 = 7'h63 == io_i_rename_table_3 ? io_i_pregs_99 : _GEN_482; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_484 = 7'h64 == io_i_rename_table_3 ? io_i_pregs_100 : _GEN_483; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_485 = 7'h65 == io_i_rename_table_3 ? io_i_pregs_101 : _GEN_484; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_486 = 7'h66 == io_i_rename_table_3 ? io_i_pregs_102 : _GEN_485; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_487 = 7'h67 == io_i_rename_table_3 ? io_i_pregs_103 : _GEN_486; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_488 = 7'h68 == io_i_rename_table_3 ? io_i_pregs_104 : _GEN_487; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_489 = 7'h69 == io_i_rename_table_3 ? io_i_pregs_105 : _GEN_488; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_490 = 7'h6a == io_i_rename_table_3 ? io_i_pregs_106 : _GEN_489; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_491 = 7'h6b == io_i_rename_table_3 ? io_i_pregs_107 : _GEN_490; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_492 = 7'h6c == io_i_rename_table_3 ? io_i_pregs_108 : _GEN_491; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_493 = 7'h6d == io_i_rename_table_3 ? io_i_pregs_109 : _GEN_492; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_494 = 7'h6e == io_i_rename_table_3 ? io_i_pregs_110 : _GEN_493; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_495 = 7'h6f == io_i_rename_table_3 ? io_i_pregs_111 : _GEN_494; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_496 = 7'h70 == io_i_rename_table_3 ? io_i_pregs_112 : _GEN_495; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_497 = 7'h71 == io_i_rename_table_3 ? io_i_pregs_113 : _GEN_496; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_498 = 7'h72 == io_i_rename_table_3 ? io_i_pregs_114 : _GEN_497; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_499 = 7'h73 == io_i_rename_table_3 ? io_i_pregs_115 : _GEN_498; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_500 = 7'h74 == io_i_rename_table_3 ? io_i_pregs_116 : _GEN_499; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_501 = 7'h75 == io_i_rename_table_3 ? io_i_pregs_117 : _GEN_500; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_502 = 7'h76 == io_i_rename_table_3 ? io_i_pregs_118 : _GEN_501; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_503 = 7'h77 == io_i_rename_table_3 ? io_i_pregs_119 : _GEN_502; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_504 = 7'h78 == io_i_rename_table_3 ? io_i_pregs_120 : _GEN_503; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_505 = 7'h79 == io_i_rename_table_3 ? io_i_pregs_121 : _GEN_504; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_506 = 7'h7a == io_i_rename_table_3 ? io_i_pregs_122 : _GEN_505; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_507 = 7'h7b == io_i_rename_table_3 ? io_i_pregs_123 : _GEN_506; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_508 = 7'h7c == io_i_rename_table_3 ? io_i_pregs_124 : _GEN_507; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_509 = 7'h7d == io_i_rename_table_3 ? io_i_pregs_125 : _GEN_508; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_510 = 7'h7e == io_i_rename_table_3 ? io_i_pregs_126 : _GEN_509; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_513 = 7'h1 == io_i_rename_table_4 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_514 = 7'h2 == io_i_rename_table_4 ? io_i_pregs_2 : _GEN_513; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_515 = 7'h3 == io_i_rename_table_4 ? io_i_pregs_3 : _GEN_514; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_516 = 7'h4 == io_i_rename_table_4 ? io_i_pregs_4 : _GEN_515; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_517 = 7'h5 == io_i_rename_table_4 ? io_i_pregs_5 : _GEN_516; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_518 = 7'h6 == io_i_rename_table_4 ? io_i_pregs_6 : _GEN_517; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_519 = 7'h7 == io_i_rename_table_4 ? io_i_pregs_7 : _GEN_518; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_520 = 7'h8 == io_i_rename_table_4 ? io_i_pregs_8 : _GEN_519; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_521 = 7'h9 == io_i_rename_table_4 ? io_i_pregs_9 : _GEN_520; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_522 = 7'ha == io_i_rename_table_4 ? io_i_pregs_10 : _GEN_521; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_523 = 7'hb == io_i_rename_table_4 ? io_i_pregs_11 : _GEN_522; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_524 = 7'hc == io_i_rename_table_4 ? io_i_pregs_12 : _GEN_523; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_525 = 7'hd == io_i_rename_table_4 ? io_i_pregs_13 : _GEN_524; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_526 = 7'he == io_i_rename_table_4 ? io_i_pregs_14 : _GEN_525; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_527 = 7'hf == io_i_rename_table_4 ? io_i_pregs_15 : _GEN_526; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_528 = 7'h10 == io_i_rename_table_4 ? io_i_pregs_16 : _GEN_527; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_529 = 7'h11 == io_i_rename_table_4 ? io_i_pregs_17 : _GEN_528; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_530 = 7'h12 == io_i_rename_table_4 ? io_i_pregs_18 : _GEN_529; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_531 = 7'h13 == io_i_rename_table_4 ? io_i_pregs_19 : _GEN_530; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_532 = 7'h14 == io_i_rename_table_4 ? io_i_pregs_20 : _GEN_531; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_533 = 7'h15 == io_i_rename_table_4 ? io_i_pregs_21 : _GEN_532; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_534 = 7'h16 == io_i_rename_table_4 ? io_i_pregs_22 : _GEN_533; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_535 = 7'h17 == io_i_rename_table_4 ? io_i_pregs_23 : _GEN_534; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_536 = 7'h18 == io_i_rename_table_4 ? io_i_pregs_24 : _GEN_535; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_537 = 7'h19 == io_i_rename_table_4 ? io_i_pregs_25 : _GEN_536; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_538 = 7'h1a == io_i_rename_table_4 ? io_i_pregs_26 : _GEN_537; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_539 = 7'h1b == io_i_rename_table_4 ? io_i_pregs_27 : _GEN_538; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_540 = 7'h1c == io_i_rename_table_4 ? io_i_pregs_28 : _GEN_539; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_541 = 7'h1d == io_i_rename_table_4 ? io_i_pregs_29 : _GEN_540; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_542 = 7'h1e == io_i_rename_table_4 ? io_i_pregs_30 : _GEN_541; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_543 = 7'h1f == io_i_rename_table_4 ? io_i_pregs_31 : _GEN_542; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_544 = 7'h20 == io_i_rename_table_4 ? io_i_pregs_32 : _GEN_543; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_545 = 7'h21 == io_i_rename_table_4 ? io_i_pregs_33 : _GEN_544; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_546 = 7'h22 == io_i_rename_table_4 ? io_i_pregs_34 : _GEN_545; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_547 = 7'h23 == io_i_rename_table_4 ? io_i_pregs_35 : _GEN_546; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_548 = 7'h24 == io_i_rename_table_4 ? io_i_pregs_36 : _GEN_547; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_549 = 7'h25 == io_i_rename_table_4 ? io_i_pregs_37 : _GEN_548; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_550 = 7'h26 == io_i_rename_table_4 ? io_i_pregs_38 : _GEN_549; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_551 = 7'h27 == io_i_rename_table_4 ? io_i_pregs_39 : _GEN_550; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_552 = 7'h28 == io_i_rename_table_4 ? io_i_pregs_40 : _GEN_551; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_553 = 7'h29 == io_i_rename_table_4 ? io_i_pregs_41 : _GEN_552; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_554 = 7'h2a == io_i_rename_table_4 ? io_i_pregs_42 : _GEN_553; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_555 = 7'h2b == io_i_rename_table_4 ? io_i_pregs_43 : _GEN_554; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_556 = 7'h2c == io_i_rename_table_4 ? io_i_pregs_44 : _GEN_555; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_557 = 7'h2d == io_i_rename_table_4 ? io_i_pregs_45 : _GEN_556; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_558 = 7'h2e == io_i_rename_table_4 ? io_i_pregs_46 : _GEN_557; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_559 = 7'h2f == io_i_rename_table_4 ? io_i_pregs_47 : _GEN_558; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_560 = 7'h30 == io_i_rename_table_4 ? io_i_pregs_48 : _GEN_559; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_561 = 7'h31 == io_i_rename_table_4 ? io_i_pregs_49 : _GEN_560; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_562 = 7'h32 == io_i_rename_table_4 ? io_i_pregs_50 : _GEN_561; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_563 = 7'h33 == io_i_rename_table_4 ? io_i_pregs_51 : _GEN_562; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_564 = 7'h34 == io_i_rename_table_4 ? io_i_pregs_52 : _GEN_563; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_565 = 7'h35 == io_i_rename_table_4 ? io_i_pregs_53 : _GEN_564; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_566 = 7'h36 == io_i_rename_table_4 ? io_i_pregs_54 : _GEN_565; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_567 = 7'h37 == io_i_rename_table_4 ? io_i_pregs_55 : _GEN_566; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_568 = 7'h38 == io_i_rename_table_4 ? io_i_pregs_56 : _GEN_567; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_569 = 7'h39 == io_i_rename_table_4 ? io_i_pregs_57 : _GEN_568; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_570 = 7'h3a == io_i_rename_table_4 ? io_i_pregs_58 : _GEN_569; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_571 = 7'h3b == io_i_rename_table_4 ? io_i_pregs_59 : _GEN_570; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_572 = 7'h3c == io_i_rename_table_4 ? io_i_pregs_60 : _GEN_571; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_573 = 7'h3d == io_i_rename_table_4 ? io_i_pregs_61 : _GEN_572; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_574 = 7'h3e == io_i_rename_table_4 ? io_i_pregs_62 : _GEN_573; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_575 = 7'h3f == io_i_rename_table_4 ? io_i_pregs_63 : _GEN_574; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_576 = 7'h40 == io_i_rename_table_4 ? io_i_pregs_64 : _GEN_575; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_577 = 7'h41 == io_i_rename_table_4 ? io_i_pregs_65 : _GEN_576; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_578 = 7'h42 == io_i_rename_table_4 ? io_i_pregs_66 : _GEN_577; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_579 = 7'h43 == io_i_rename_table_4 ? io_i_pregs_67 : _GEN_578; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_580 = 7'h44 == io_i_rename_table_4 ? io_i_pregs_68 : _GEN_579; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_581 = 7'h45 == io_i_rename_table_4 ? io_i_pregs_69 : _GEN_580; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_582 = 7'h46 == io_i_rename_table_4 ? io_i_pregs_70 : _GEN_581; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_583 = 7'h47 == io_i_rename_table_4 ? io_i_pregs_71 : _GEN_582; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_584 = 7'h48 == io_i_rename_table_4 ? io_i_pregs_72 : _GEN_583; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_585 = 7'h49 == io_i_rename_table_4 ? io_i_pregs_73 : _GEN_584; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_586 = 7'h4a == io_i_rename_table_4 ? io_i_pregs_74 : _GEN_585; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_587 = 7'h4b == io_i_rename_table_4 ? io_i_pregs_75 : _GEN_586; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_588 = 7'h4c == io_i_rename_table_4 ? io_i_pregs_76 : _GEN_587; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_589 = 7'h4d == io_i_rename_table_4 ? io_i_pregs_77 : _GEN_588; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_590 = 7'h4e == io_i_rename_table_4 ? io_i_pregs_78 : _GEN_589; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_591 = 7'h4f == io_i_rename_table_4 ? io_i_pregs_79 : _GEN_590; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_592 = 7'h50 == io_i_rename_table_4 ? io_i_pregs_80 : _GEN_591; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_593 = 7'h51 == io_i_rename_table_4 ? io_i_pregs_81 : _GEN_592; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_594 = 7'h52 == io_i_rename_table_4 ? io_i_pregs_82 : _GEN_593; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_595 = 7'h53 == io_i_rename_table_4 ? io_i_pregs_83 : _GEN_594; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_596 = 7'h54 == io_i_rename_table_4 ? io_i_pregs_84 : _GEN_595; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_597 = 7'h55 == io_i_rename_table_4 ? io_i_pregs_85 : _GEN_596; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_598 = 7'h56 == io_i_rename_table_4 ? io_i_pregs_86 : _GEN_597; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_599 = 7'h57 == io_i_rename_table_4 ? io_i_pregs_87 : _GEN_598; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_600 = 7'h58 == io_i_rename_table_4 ? io_i_pregs_88 : _GEN_599; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_601 = 7'h59 == io_i_rename_table_4 ? io_i_pregs_89 : _GEN_600; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_602 = 7'h5a == io_i_rename_table_4 ? io_i_pregs_90 : _GEN_601; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_603 = 7'h5b == io_i_rename_table_4 ? io_i_pregs_91 : _GEN_602; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_604 = 7'h5c == io_i_rename_table_4 ? io_i_pregs_92 : _GEN_603; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_605 = 7'h5d == io_i_rename_table_4 ? io_i_pregs_93 : _GEN_604; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_606 = 7'h5e == io_i_rename_table_4 ? io_i_pregs_94 : _GEN_605; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_607 = 7'h5f == io_i_rename_table_4 ? io_i_pregs_95 : _GEN_606; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_608 = 7'h60 == io_i_rename_table_4 ? io_i_pregs_96 : _GEN_607; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_609 = 7'h61 == io_i_rename_table_4 ? io_i_pregs_97 : _GEN_608; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_610 = 7'h62 == io_i_rename_table_4 ? io_i_pregs_98 : _GEN_609; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_611 = 7'h63 == io_i_rename_table_4 ? io_i_pregs_99 : _GEN_610; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_612 = 7'h64 == io_i_rename_table_4 ? io_i_pregs_100 : _GEN_611; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_613 = 7'h65 == io_i_rename_table_4 ? io_i_pregs_101 : _GEN_612; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_614 = 7'h66 == io_i_rename_table_4 ? io_i_pregs_102 : _GEN_613; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_615 = 7'h67 == io_i_rename_table_4 ? io_i_pregs_103 : _GEN_614; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_616 = 7'h68 == io_i_rename_table_4 ? io_i_pregs_104 : _GEN_615; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_617 = 7'h69 == io_i_rename_table_4 ? io_i_pregs_105 : _GEN_616; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_618 = 7'h6a == io_i_rename_table_4 ? io_i_pregs_106 : _GEN_617; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_619 = 7'h6b == io_i_rename_table_4 ? io_i_pregs_107 : _GEN_618; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_620 = 7'h6c == io_i_rename_table_4 ? io_i_pregs_108 : _GEN_619; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_621 = 7'h6d == io_i_rename_table_4 ? io_i_pregs_109 : _GEN_620; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_622 = 7'h6e == io_i_rename_table_4 ? io_i_pregs_110 : _GEN_621; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_623 = 7'h6f == io_i_rename_table_4 ? io_i_pregs_111 : _GEN_622; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_624 = 7'h70 == io_i_rename_table_4 ? io_i_pregs_112 : _GEN_623; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_625 = 7'h71 == io_i_rename_table_4 ? io_i_pregs_113 : _GEN_624; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_626 = 7'h72 == io_i_rename_table_4 ? io_i_pregs_114 : _GEN_625; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_627 = 7'h73 == io_i_rename_table_4 ? io_i_pregs_115 : _GEN_626; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_628 = 7'h74 == io_i_rename_table_4 ? io_i_pregs_116 : _GEN_627; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_629 = 7'h75 == io_i_rename_table_4 ? io_i_pregs_117 : _GEN_628; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_630 = 7'h76 == io_i_rename_table_4 ? io_i_pregs_118 : _GEN_629; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_631 = 7'h77 == io_i_rename_table_4 ? io_i_pregs_119 : _GEN_630; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_632 = 7'h78 == io_i_rename_table_4 ? io_i_pregs_120 : _GEN_631; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_633 = 7'h79 == io_i_rename_table_4 ? io_i_pregs_121 : _GEN_632; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_634 = 7'h7a == io_i_rename_table_4 ? io_i_pregs_122 : _GEN_633; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_635 = 7'h7b == io_i_rename_table_4 ? io_i_pregs_123 : _GEN_634; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_636 = 7'h7c == io_i_rename_table_4 ? io_i_pregs_124 : _GEN_635; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_637 = 7'h7d == io_i_rename_table_4 ? io_i_pregs_125 : _GEN_636; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_638 = 7'h7e == io_i_rename_table_4 ? io_i_pregs_126 : _GEN_637; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_641 = 7'h1 == io_i_rename_table_5 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_642 = 7'h2 == io_i_rename_table_5 ? io_i_pregs_2 : _GEN_641; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_643 = 7'h3 == io_i_rename_table_5 ? io_i_pregs_3 : _GEN_642; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_644 = 7'h4 == io_i_rename_table_5 ? io_i_pregs_4 : _GEN_643; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_645 = 7'h5 == io_i_rename_table_5 ? io_i_pregs_5 : _GEN_644; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_646 = 7'h6 == io_i_rename_table_5 ? io_i_pregs_6 : _GEN_645; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_647 = 7'h7 == io_i_rename_table_5 ? io_i_pregs_7 : _GEN_646; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_648 = 7'h8 == io_i_rename_table_5 ? io_i_pregs_8 : _GEN_647; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_649 = 7'h9 == io_i_rename_table_5 ? io_i_pregs_9 : _GEN_648; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_650 = 7'ha == io_i_rename_table_5 ? io_i_pregs_10 : _GEN_649; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_651 = 7'hb == io_i_rename_table_5 ? io_i_pregs_11 : _GEN_650; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_652 = 7'hc == io_i_rename_table_5 ? io_i_pregs_12 : _GEN_651; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_653 = 7'hd == io_i_rename_table_5 ? io_i_pregs_13 : _GEN_652; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_654 = 7'he == io_i_rename_table_5 ? io_i_pregs_14 : _GEN_653; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_655 = 7'hf == io_i_rename_table_5 ? io_i_pregs_15 : _GEN_654; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_656 = 7'h10 == io_i_rename_table_5 ? io_i_pregs_16 : _GEN_655; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_657 = 7'h11 == io_i_rename_table_5 ? io_i_pregs_17 : _GEN_656; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_658 = 7'h12 == io_i_rename_table_5 ? io_i_pregs_18 : _GEN_657; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_659 = 7'h13 == io_i_rename_table_5 ? io_i_pregs_19 : _GEN_658; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_660 = 7'h14 == io_i_rename_table_5 ? io_i_pregs_20 : _GEN_659; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_661 = 7'h15 == io_i_rename_table_5 ? io_i_pregs_21 : _GEN_660; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_662 = 7'h16 == io_i_rename_table_5 ? io_i_pregs_22 : _GEN_661; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_663 = 7'h17 == io_i_rename_table_5 ? io_i_pregs_23 : _GEN_662; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_664 = 7'h18 == io_i_rename_table_5 ? io_i_pregs_24 : _GEN_663; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_665 = 7'h19 == io_i_rename_table_5 ? io_i_pregs_25 : _GEN_664; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_666 = 7'h1a == io_i_rename_table_5 ? io_i_pregs_26 : _GEN_665; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_667 = 7'h1b == io_i_rename_table_5 ? io_i_pregs_27 : _GEN_666; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_668 = 7'h1c == io_i_rename_table_5 ? io_i_pregs_28 : _GEN_667; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_669 = 7'h1d == io_i_rename_table_5 ? io_i_pregs_29 : _GEN_668; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_670 = 7'h1e == io_i_rename_table_5 ? io_i_pregs_30 : _GEN_669; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_671 = 7'h1f == io_i_rename_table_5 ? io_i_pregs_31 : _GEN_670; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_672 = 7'h20 == io_i_rename_table_5 ? io_i_pregs_32 : _GEN_671; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_673 = 7'h21 == io_i_rename_table_5 ? io_i_pregs_33 : _GEN_672; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_674 = 7'h22 == io_i_rename_table_5 ? io_i_pregs_34 : _GEN_673; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_675 = 7'h23 == io_i_rename_table_5 ? io_i_pregs_35 : _GEN_674; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_676 = 7'h24 == io_i_rename_table_5 ? io_i_pregs_36 : _GEN_675; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_677 = 7'h25 == io_i_rename_table_5 ? io_i_pregs_37 : _GEN_676; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_678 = 7'h26 == io_i_rename_table_5 ? io_i_pregs_38 : _GEN_677; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_679 = 7'h27 == io_i_rename_table_5 ? io_i_pregs_39 : _GEN_678; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_680 = 7'h28 == io_i_rename_table_5 ? io_i_pregs_40 : _GEN_679; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_681 = 7'h29 == io_i_rename_table_5 ? io_i_pregs_41 : _GEN_680; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_682 = 7'h2a == io_i_rename_table_5 ? io_i_pregs_42 : _GEN_681; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_683 = 7'h2b == io_i_rename_table_5 ? io_i_pregs_43 : _GEN_682; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_684 = 7'h2c == io_i_rename_table_5 ? io_i_pregs_44 : _GEN_683; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_685 = 7'h2d == io_i_rename_table_5 ? io_i_pregs_45 : _GEN_684; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_686 = 7'h2e == io_i_rename_table_5 ? io_i_pregs_46 : _GEN_685; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_687 = 7'h2f == io_i_rename_table_5 ? io_i_pregs_47 : _GEN_686; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_688 = 7'h30 == io_i_rename_table_5 ? io_i_pregs_48 : _GEN_687; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_689 = 7'h31 == io_i_rename_table_5 ? io_i_pregs_49 : _GEN_688; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_690 = 7'h32 == io_i_rename_table_5 ? io_i_pregs_50 : _GEN_689; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_691 = 7'h33 == io_i_rename_table_5 ? io_i_pregs_51 : _GEN_690; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_692 = 7'h34 == io_i_rename_table_5 ? io_i_pregs_52 : _GEN_691; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_693 = 7'h35 == io_i_rename_table_5 ? io_i_pregs_53 : _GEN_692; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_694 = 7'h36 == io_i_rename_table_5 ? io_i_pregs_54 : _GEN_693; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_695 = 7'h37 == io_i_rename_table_5 ? io_i_pregs_55 : _GEN_694; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_696 = 7'h38 == io_i_rename_table_5 ? io_i_pregs_56 : _GEN_695; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_697 = 7'h39 == io_i_rename_table_5 ? io_i_pregs_57 : _GEN_696; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_698 = 7'h3a == io_i_rename_table_5 ? io_i_pregs_58 : _GEN_697; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_699 = 7'h3b == io_i_rename_table_5 ? io_i_pregs_59 : _GEN_698; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_700 = 7'h3c == io_i_rename_table_5 ? io_i_pregs_60 : _GEN_699; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_701 = 7'h3d == io_i_rename_table_5 ? io_i_pregs_61 : _GEN_700; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_702 = 7'h3e == io_i_rename_table_5 ? io_i_pregs_62 : _GEN_701; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_703 = 7'h3f == io_i_rename_table_5 ? io_i_pregs_63 : _GEN_702; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_704 = 7'h40 == io_i_rename_table_5 ? io_i_pregs_64 : _GEN_703; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_705 = 7'h41 == io_i_rename_table_5 ? io_i_pregs_65 : _GEN_704; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_706 = 7'h42 == io_i_rename_table_5 ? io_i_pregs_66 : _GEN_705; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_707 = 7'h43 == io_i_rename_table_5 ? io_i_pregs_67 : _GEN_706; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_708 = 7'h44 == io_i_rename_table_5 ? io_i_pregs_68 : _GEN_707; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_709 = 7'h45 == io_i_rename_table_5 ? io_i_pregs_69 : _GEN_708; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_710 = 7'h46 == io_i_rename_table_5 ? io_i_pregs_70 : _GEN_709; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_711 = 7'h47 == io_i_rename_table_5 ? io_i_pregs_71 : _GEN_710; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_712 = 7'h48 == io_i_rename_table_5 ? io_i_pregs_72 : _GEN_711; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_713 = 7'h49 == io_i_rename_table_5 ? io_i_pregs_73 : _GEN_712; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_714 = 7'h4a == io_i_rename_table_5 ? io_i_pregs_74 : _GEN_713; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_715 = 7'h4b == io_i_rename_table_5 ? io_i_pregs_75 : _GEN_714; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_716 = 7'h4c == io_i_rename_table_5 ? io_i_pregs_76 : _GEN_715; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_717 = 7'h4d == io_i_rename_table_5 ? io_i_pregs_77 : _GEN_716; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_718 = 7'h4e == io_i_rename_table_5 ? io_i_pregs_78 : _GEN_717; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_719 = 7'h4f == io_i_rename_table_5 ? io_i_pregs_79 : _GEN_718; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_720 = 7'h50 == io_i_rename_table_5 ? io_i_pregs_80 : _GEN_719; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_721 = 7'h51 == io_i_rename_table_5 ? io_i_pregs_81 : _GEN_720; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_722 = 7'h52 == io_i_rename_table_5 ? io_i_pregs_82 : _GEN_721; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_723 = 7'h53 == io_i_rename_table_5 ? io_i_pregs_83 : _GEN_722; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_724 = 7'h54 == io_i_rename_table_5 ? io_i_pregs_84 : _GEN_723; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_725 = 7'h55 == io_i_rename_table_5 ? io_i_pregs_85 : _GEN_724; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_726 = 7'h56 == io_i_rename_table_5 ? io_i_pregs_86 : _GEN_725; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_727 = 7'h57 == io_i_rename_table_5 ? io_i_pregs_87 : _GEN_726; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_728 = 7'h58 == io_i_rename_table_5 ? io_i_pregs_88 : _GEN_727; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_729 = 7'h59 == io_i_rename_table_5 ? io_i_pregs_89 : _GEN_728; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_730 = 7'h5a == io_i_rename_table_5 ? io_i_pregs_90 : _GEN_729; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_731 = 7'h5b == io_i_rename_table_5 ? io_i_pregs_91 : _GEN_730; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_732 = 7'h5c == io_i_rename_table_5 ? io_i_pregs_92 : _GEN_731; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_733 = 7'h5d == io_i_rename_table_5 ? io_i_pregs_93 : _GEN_732; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_734 = 7'h5e == io_i_rename_table_5 ? io_i_pregs_94 : _GEN_733; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_735 = 7'h5f == io_i_rename_table_5 ? io_i_pregs_95 : _GEN_734; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_736 = 7'h60 == io_i_rename_table_5 ? io_i_pregs_96 : _GEN_735; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_737 = 7'h61 == io_i_rename_table_5 ? io_i_pregs_97 : _GEN_736; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_738 = 7'h62 == io_i_rename_table_5 ? io_i_pregs_98 : _GEN_737; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_739 = 7'h63 == io_i_rename_table_5 ? io_i_pregs_99 : _GEN_738; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_740 = 7'h64 == io_i_rename_table_5 ? io_i_pregs_100 : _GEN_739; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_741 = 7'h65 == io_i_rename_table_5 ? io_i_pregs_101 : _GEN_740; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_742 = 7'h66 == io_i_rename_table_5 ? io_i_pregs_102 : _GEN_741; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_743 = 7'h67 == io_i_rename_table_5 ? io_i_pregs_103 : _GEN_742; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_744 = 7'h68 == io_i_rename_table_5 ? io_i_pregs_104 : _GEN_743; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_745 = 7'h69 == io_i_rename_table_5 ? io_i_pregs_105 : _GEN_744; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_746 = 7'h6a == io_i_rename_table_5 ? io_i_pregs_106 : _GEN_745; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_747 = 7'h6b == io_i_rename_table_5 ? io_i_pregs_107 : _GEN_746; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_748 = 7'h6c == io_i_rename_table_5 ? io_i_pregs_108 : _GEN_747; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_749 = 7'h6d == io_i_rename_table_5 ? io_i_pregs_109 : _GEN_748; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_750 = 7'h6e == io_i_rename_table_5 ? io_i_pregs_110 : _GEN_749; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_751 = 7'h6f == io_i_rename_table_5 ? io_i_pregs_111 : _GEN_750; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_752 = 7'h70 == io_i_rename_table_5 ? io_i_pregs_112 : _GEN_751; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_753 = 7'h71 == io_i_rename_table_5 ? io_i_pregs_113 : _GEN_752; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_754 = 7'h72 == io_i_rename_table_5 ? io_i_pregs_114 : _GEN_753; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_755 = 7'h73 == io_i_rename_table_5 ? io_i_pregs_115 : _GEN_754; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_756 = 7'h74 == io_i_rename_table_5 ? io_i_pregs_116 : _GEN_755; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_757 = 7'h75 == io_i_rename_table_5 ? io_i_pregs_117 : _GEN_756; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_758 = 7'h76 == io_i_rename_table_5 ? io_i_pregs_118 : _GEN_757; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_759 = 7'h77 == io_i_rename_table_5 ? io_i_pregs_119 : _GEN_758; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_760 = 7'h78 == io_i_rename_table_5 ? io_i_pregs_120 : _GEN_759; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_761 = 7'h79 == io_i_rename_table_5 ? io_i_pregs_121 : _GEN_760; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_762 = 7'h7a == io_i_rename_table_5 ? io_i_pregs_122 : _GEN_761; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_763 = 7'h7b == io_i_rename_table_5 ? io_i_pregs_123 : _GEN_762; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_764 = 7'h7c == io_i_rename_table_5 ? io_i_pregs_124 : _GEN_763; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_765 = 7'h7d == io_i_rename_table_5 ? io_i_pregs_125 : _GEN_764; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_766 = 7'h7e == io_i_rename_table_5 ? io_i_pregs_126 : _GEN_765; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_769 = 7'h1 == io_i_rename_table_6 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_770 = 7'h2 == io_i_rename_table_6 ? io_i_pregs_2 : _GEN_769; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_771 = 7'h3 == io_i_rename_table_6 ? io_i_pregs_3 : _GEN_770; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_772 = 7'h4 == io_i_rename_table_6 ? io_i_pregs_4 : _GEN_771; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_773 = 7'h5 == io_i_rename_table_6 ? io_i_pregs_5 : _GEN_772; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_774 = 7'h6 == io_i_rename_table_6 ? io_i_pregs_6 : _GEN_773; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_775 = 7'h7 == io_i_rename_table_6 ? io_i_pregs_7 : _GEN_774; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_776 = 7'h8 == io_i_rename_table_6 ? io_i_pregs_8 : _GEN_775; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_777 = 7'h9 == io_i_rename_table_6 ? io_i_pregs_9 : _GEN_776; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_778 = 7'ha == io_i_rename_table_6 ? io_i_pregs_10 : _GEN_777; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_779 = 7'hb == io_i_rename_table_6 ? io_i_pregs_11 : _GEN_778; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_780 = 7'hc == io_i_rename_table_6 ? io_i_pregs_12 : _GEN_779; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_781 = 7'hd == io_i_rename_table_6 ? io_i_pregs_13 : _GEN_780; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_782 = 7'he == io_i_rename_table_6 ? io_i_pregs_14 : _GEN_781; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_783 = 7'hf == io_i_rename_table_6 ? io_i_pregs_15 : _GEN_782; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_784 = 7'h10 == io_i_rename_table_6 ? io_i_pregs_16 : _GEN_783; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_785 = 7'h11 == io_i_rename_table_6 ? io_i_pregs_17 : _GEN_784; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_786 = 7'h12 == io_i_rename_table_6 ? io_i_pregs_18 : _GEN_785; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_787 = 7'h13 == io_i_rename_table_6 ? io_i_pregs_19 : _GEN_786; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_788 = 7'h14 == io_i_rename_table_6 ? io_i_pregs_20 : _GEN_787; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_789 = 7'h15 == io_i_rename_table_6 ? io_i_pregs_21 : _GEN_788; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_790 = 7'h16 == io_i_rename_table_6 ? io_i_pregs_22 : _GEN_789; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_791 = 7'h17 == io_i_rename_table_6 ? io_i_pregs_23 : _GEN_790; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_792 = 7'h18 == io_i_rename_table_6 ? io_i_pregs_24 : _GEN_791; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_793 = 7'h19 == io_i_rename_table_6 ? io_i_pregs_25 : _GEN_792; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_794 = 7'h1a == io_i_rename_table_6 ? io_i_pregs_26 : _GEN_793; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_795 = 7'h1b == io_i_rename_table_6 ? io_i_pregs_27 : _GEN_794; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_796 = 7'h1c == io_i_rename_table_6 ? io_i_pregs_28 : _GEN_795; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_797 = 7'h1d == io_i_rename_table_6 ? io_i_pregs_29 : _GEN_796; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_798 = 7'h1e == io_i_rename_table_6 ? io_i_pregs_30 : _GEN_797; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_799 = 7'h1f == io_i_rename_table_6 ? io_i_pregs_31 : _GEN_798; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_800 = 7'h20 == io_i_rename_table_6 ? io_i_pregs_32 : _GEN_799; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_801 = 7'h21 == io_i_rename_table_6 ? io_i_pregs_33 : _GEN_800; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_802 = 7'h22 == io_i_rename_table_6 ? io_i_pregs_34 : _GEN_801; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_803 = 7'h23 == io_i_rename_table_6 ? io_i_pregs_35 : _GEN_802; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_804 = 7'h24 == io_i_rename_table_6 ? io_i_pregs_36 : _GEN_803; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_805 = 7'h25 == io_i_rename_table_6 ? io_i_pregs_37 : _GEN_804; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_806 = 7'h26 == io_i_rename_table_6 ? io_i_pregs_38 : _GEN_805; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_807 = 7'h27 == io_i_rename_table_6 ? io_i_pregs_39 : _GEN_806; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_808 = 7'h28 == io_i_rename_table_6 ? io_i_pregs_40 : _GEN_807; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_809 = 7'h29 == io_i_rename_table_6 ? io_i_pregs_41 : _GEN_808; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_810 = 7'h2a == io_i_rename_table_6 ? io_i_pregs_42 : _GEN_809; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_811 = 7'h2b == io_i_rename_table_6 ? io_i_pregs_43 : _GEN_810; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_812 = 7'h2c == io_i_rename_table_6 ? io_i_pregs_44 : _GEN_811; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_813 = 7'h2d == io_i_rename_table_6 ? io_i_pregs_45 : _GEN_812; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_814 = 7'h2e == io_i_rename_table_6 ? io_i_pregs_46 : _GEN_813; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_815 = 7'h2f == io_i_rename_table_6 ? io_i_pregs_47 : _GEN_814; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_816 = 7'h30 == io_i_rename_table_6 ? io_i_pregs_48 : _GEN_815; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_817 = 7'h31 == io_i_rename_table_6 ? io_i_pregs_49 : _GEN_816; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_818 = 7'h32 == io_i_rename_table_6 ? io_i_pregs_50 : _GEN_817; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_819 = 7'h33 == io_i_rename_table_6 ? io_i_pregs_51 : _GEN_818; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_820 = 7'h34 == io_i_rename_table_6 ? io_i_pregs_52 : _GEN_819; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_821 = 7'h35 == io_i_rename_table_6 ? io_i_pregs_53 : _GEN_820; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_822 = 7'h36 == io_i_rename_table_6 ? io_i_pregs_54 : _GEN_821; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_823 = 7'h37 == io_i_rename_table_6 ? io_i_pregs_55 : _GEN_822; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_824 = 7'h38 == io_i_rename_table_6 ? io_i_pregs_56 : _GEN_823; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_825 = 7'h39 == io_i_rename_table_6 ? io_i_pregs_57 : _GEN_824; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_826 = 7'h3a == io_i_rename_table_6 ? io_i_pregs_58 : _GEN_825; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_827 = 7'h3b == io_i_rename_table_6 ? io_i_pregs_59 : _GEN_826; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_828 = 7'h3c == io_i_rename_table_6 ? io_i_pregs_60 : _GEN_827; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_829 = 7'h3d == io_i_rename_table_6 ? io_i_pregs_61 : _GEN_828; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_830 = 7'h3e == io_i_rename_table_6 ? io_i_pregs_62 : _GEN_829; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_831 = 7'h3f == io_i_rename_table_6 ? io_i_pregs_63 : _GEN_830; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_832 = 7'h40 == io_i_rename_table_6 ? io_i_pregs_64 : _GEN_831; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_833 = 7'h41 == io_i_rename_table_6 ? io_i_pregs_65 : _GEN_832; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_834 = 7'h42 == io_i_rename_table_6 ? io_i_pregs_66 : _GEN_833; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_835 = 7'h43 == io_i_rename_table_6 ? io_i_pregs_67 : _GEN_834; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_836 = 7'h44 == io_i_rename_table_6 ? io_i_pregs_68 : _GEN_835; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_837 = 7'h45 == io_i_rename_table_6 ? io_i_pregs_69 : _GEN_836; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_838 = 7'h46 == io_i_rename_table_6 ? io_i_pregs_70 : _GEN_837; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_839 = 7'h47 == io_i_rename_table_6 ? io_i_pregs_71 : _GEN_838; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_840 = 7'h48 == io_i_rename_table_6 ? io_i_pregs_72 : _GEN_839; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_841 = 7'h49 == io_i_rename_table_6 ? io_i_pregs_73 : _GEN_840; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_842 = 7'h4a == io_i_rename_table_6 ? io_i_pregs_74 : _GEN_841; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_843 = 7'h4b == io_i_rename_table_6 ? io_i_pregs_75 : _GEN_842; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_844 = 7'h4c == io_i_rename_table_6 ? io_i_pregs_76 : _GEN_843; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_845 = 7'h4d == io_i_rename_table_6 ? io_i_pregs_77 : _GEN_844; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_846 = 7'h4e == io_i_rename_table_6 ? io_i_pregs_78 : _GEN_845; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_847 = 7'h4f == io_i_rename_table_6 ? io_i_pregs_79 : _GEN_846; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_848 = 7'h50 == io_i_rename_table_6 ? io_i_pregs_80 : _GEN_847; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_849 = 7'h51 == io_i_rename_table_6 ? io_i_pregs_81 : _GEN_848; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_850 = 7'h52 == io_i_rename_table_6 ? io_i_pregs_82 : _GEN_849; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_851 = 7'h53 == io_i_rename_table_6 ? io_i_pregs_83 : _GEN_850; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_852 = 7'h54 == io_i_rename_table_6 ? io_i_pregs_84 : _GEN_851; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_853 = 7'h55 == io_i_rename_table_6 ? io_i_pregs_85 : _GEN_852; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_854 = 7'h56 == io_i_rename_table_6 ? io_i_pregs_86 : _GEN_853; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_855 = 7'h57 == io_i_rename_table_6 ? io_i_pregs_87 : _GEN_854; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_856 = 7'h58 == io_i_rename_table_6 ? io_i_pregs_88 : _GEN_855; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_857 = 7'h59 == io_i_rename_table_6 ? io_i_pregs_89 : _GEN_856; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_858 = 7'h5a == io_i_rename_table_6 ? io_i_pregs_90 : _GEN_857; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_859 = 7'h5b == io_i_rename_table_6 ? io_i_pregs_91 : _GEN_858; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_860 = 7'h5c == io_i_rename_table_6 ? io_i_pregs_92 : _GEN_859; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_861 = 7'h5d == io_i_rename_table_6 ? io_i_pregs_93 : _GEN_860; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_862 = 7'h5e == io_i_rename_table_6 ? io_i_pregs_94 : _GEN_861; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_863 = 7'h5f == io_i_rename_table_6 ? io_i_pregs_95 : _GEN_862; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_864 = 7'h60 == io_i_rename_table_6 ? io_i_pregs_96 : _GEN_863; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_865 = 7'h61 == io_i_rename_table_6 ? io_i_pregs_97 : _GEN_864; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_866 = 7'h62 == io_i_rename_table_6 ? io_i_pregs_98 : _GEN_865; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_867 = 7'h63 == io_i_rename_table_6 ? io_i_pregs_99 : _GEN_866; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_868 = 7'h64 == io_i_rename_table_6 ? io_i_pregs_100 : _GEN_867; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_869 = 7'h65 == io_i_rename_table_6 ? io_i_pregs_101 : _GEN_868; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_870 = 7'h66 == io_i_rename_table_6 ? io_i_pregs_102 : _GEN_869; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_871 = 7'h67 == io_i_rename_table_6 ? io_i_pregs_103 : _GEN_870; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_872 = 7'h68 == io_i_rename_table_6 ? io_i_pregs_104 : _GEN_871; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_873 = 7'h69 == io_i_rename_table_6 ? io_i_pregs_105 : _GEN_872; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_874 = 7'h6a == io_i_rename_table_6 ? io_i_pregs_106 : _GEN_873; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_875 = 7'h6b == io_i_rename_table_6 ? io_i_pregs_107 : _GEN_874; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_876 = 7'h6c == io_i_rename_table_6 ? io_i_pregs_108 : _GEN_875; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_877 = 7'h6d == io_i_rename_table_6 ? io_i_pregs_109 : _GEN_876; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_878 = 7'h6e == io_i_rename_table_6 ? io_i_pregs_110 : _GEN_877; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_879 = 7'h6f == io_i_rename_table_6 ? io_i_pregs_111 : _GEN_878; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_880 = 7'h70 == io_i_rename_table_6 ? io_i_pregs_112 : _GEN_879; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_881 = 7'h71 == io_i_rename_table_6 ? io_i_pregs_113 : _GEN_880; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_882 = 7'h72 == io_i_rename_table_6 ? io_i_pregs_114 : _GEN_881; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_883 = 7'h73 == io_i_rename_table_6 ? io_i_pregs_115 : _GEN_882; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_884 = 7'h74 == io_i_rename_table_6 ? io_i_pregs_116 : _GEN_883; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_885 = 7'h75 == io_i_rename_table_6 ? io_i_pregs_117 : _GEN_884; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_886 = 7'h76 == io_i_rename_table_6 ? io_i_pregs_118 : _GEN_885; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_887 = 7'h77 == io_i_rename_table_6 ? io_i_pregs_119 : _GEN_886; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_888 = 7'h78 == io_i_rename_table_6 ? io_i_pregs_120 : _GEN_887; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_889 = 7'h79 == io_i_rename_table_6 ? io_i_pregs_121 : _GEN_888; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_890 = 7'h7a == io_i_rename_table_6 ? io_i_pregs_122 : _GEN_889; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_891 = 7'h7b == io_i_rename_table_6 ? io_i_pregs_123 : _GEN_890; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_892 = 7'h7c == io_i_rename_table_6 ? io_i_pregs_124 : _GEN_891; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_893 = 7'h7d == io_i_rename_table_6 ? io_i_pregs_125 : _GEN_892; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_894 = 7'h7e == io_i_rename_table_6 ? io_i_pregs_126 : _GEN_893; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_897 = 7'h1 == io_i_rename_table_7 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_898 = 7'h2 == io_i_rename_table_7 ? io_i_pregs_2 : _GEN_897; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_899 = 7'h3 == io_i_rename_table_7 ? io_i_pregs_3 : _GEN_898; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_900 = 7'h4 == io_i_rename_table_7 ? io_i_pregs_4 : _GEN_899; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_901 = 7'h5 == io_i_rename_table_7 ? io_i_pregs_5 : _GEN_900; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_902 = 7'h6 == io_i_rename_table_7 ? io_i_pregs_6 : _GEN_901; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_903 = 7'h7 == io_i_rename_table_7 ? io_i_pregs_7 : _GEN_902; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_904 = 7'h8 == io_i_rename_table_7 ? io_i_pregs_8 : _GEN_903; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_905 = 7'h9 == io_i_rename_table_7 ? io_i_pregs_9 : _GEN_904; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_906 = 7'ha == io_i_rename_table_7 ? io_i_pregs_10 : _GEN_905; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_907 = 7'hb == io_i_rename_table_7 ? io_i_pregs_11 : _GEN_906; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_908 = 7'hc == io_i_rename_table_7 ? io_i_pregs_12 : _GEN_907; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_909 = 7'hd == io_i_rename_table_7 ? io_i_pregs_13 : _GEN_908; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_910 = 7'he == io_i_rename_table_7 ? io_i_pregs_14 : _GEN_909; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_911 = 7'hf == io_i_rename_table_7 ? io_i_pregs_15 : _GEN_910; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_912 = 7'h10 == io_i_rename_table_7 ? io_i_pregs_16 : _GEN_911; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_913 = 7'h11 == io_i_rename_table_7 ? io_i_pregs_17 : _GEN_912; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_914 = 7'h12 == io_i_rename_table_7 ? io_i_pregs_18 : _GEN_913; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_915 = 7'h13 == io_i_rename_table_7 ? io_i_pregs_19 : _GEN_914; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_916 = 7'h14 == io_i_rename_table_7 ? io_i_pregs_20 : _GEN_915; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_917 = 7'h15 == io_i_rename_table_7 ? io_i_pregs_21 : _GEN_916; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_918 = 7'h16 == io_i_rename_table_7 ? io_i_pregs_22 : _GEN_917; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_919 = 7'h17 == io_i_rename_table_7 ? io_i_pregs_23 : _GEN_918; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_920 = 7'h18 == io_i_rename_table_7 ? io_i_pregs_24 : _GEN_919; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_921 = 7'h19 == io_i_rename_table_7 ? io_i_pregs_25 : _GEN_920; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_922 = 7'h1a == io_i_rename_table_7 ? io_i_pregs_26 : _GEN_921; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_923 = 7'h1b == io_i_rename_table_7 ? io_i_pregs_27 : _GEN_922; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_924 = 7'h1c == io_i_rename_table_7 ? io_i_pregs_28 : _GEN_923; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_925 = 7'h1d == io_i_rename_table_7 ? io_i_pregs_29 : _GEN_924; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_926 = 7'h1e == io_i_rename_table_7 ? io_i_pregs_30 : _GEN_925; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_927 = 7'h1f == io_i_rename_table_7 ? io_i_pregs_31 : _GEN_926; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_928 = 7'h20 == io_i_rename_table_7 ? io_i_pregs_32 : _GEN_927; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_929 = 7'h21 == io_i_rename_table_7 ? io_i_pregs_33 : _GEN_928; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_930 = 7'h22 == io_i_rename_table_7 ? io_i_pregs_34 : _GEN_929; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_931 = 7'h23 == io_i_rename_table_7 ? io_i_pregs_35 : _GEN_930; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_932 = 7'h24 == io_i_rename_table_7 ? io_i_pregs_36 : _GEN_931; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_933 = 7'h25 == io_i_rename_table_7 ? io_i_pregs_37 : _GEN_932; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_934 = 7'h26 == io_i_rename_table_7 ? io_i_pregs_38 : _GEN_933; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_935 = 7'h27 == io_i_rename_table_7 ? io_i_pregs_39 : _GEN_934; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_936 = 7'h28 == io_i_rename_table_7 ? io_i_pregs_40 : _GEN_935; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_937 = 7'h29 == io_i_rename_table_7 ? io_i_pregs_41 : _GEN_936; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_938 = 7'h2a == io_i_rename_table_7 ? io_i_pregs_42 : _GEN_937; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_939 = 7'h2b == io_i_rename_table_7 ? io_i_pregs_43 : _GEN_938; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_940 = 7'h2c == io_i_rename_table_7 ? io_i_pregs_44 : _GEN_939; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_941 = 7'h2d == io_i_rename_table_7 ? io_i_pregs_45 : _GEN_940; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_942 = 7'h2e == io_i_rename_table_7 ? io_i_pregs_46 : _GEN_941; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_943 = 7'h2f == io_i_rename_table_7 ? io_i_pregs_47 : _GEN_942; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_944 = 7'h30 == io_i_rename_table_7 ? io_i_pregs_48 : _GEN_943; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_945 = 7'h31 == io_i_rename_table_7 ? io_i_pregs_49 : _GEN_944; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_946 = 7'h32 == io_i_rename_table_7 ? io_i_pregs_50 : _GEN_945; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_947 = 7'h33 == io_i_rename_table_7 ? io_i_pregs_51 : _GEN_946; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_948 = 7'h34 == io_i_rename_table_7 ? io_i_pregs_52 : _GEN_947; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_949 = 7'h35 == io_i_rename_table_7 ? io_i_pregs_53 : _GEN_948; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_950 = 7'h36 == io_i_rename_table_7 ? io_i_pregs_54 : _GEN_949; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_951 = 7'h37 == io_i_rename_table_7 ? io_i_pregs_55 : _GEN_950; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_952 = 7'h38 == io_i_rename_table_7 ? io_i_pregs_56 : _GEN_951; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_953 = 7'h39 == io_i_rename_table_7 ? io_i_pregs_57 : _GEN_952; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_954 = 7'h3a == io_i_rename_table_7 ? io_i_pregs_58 : _GEN_953; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_955 = 7'h3b == io_i_rename_table_7 ? io_i_pregs_59 : _GEN_954; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_956 = 7'h3c == io_i_rename_table_7 ? io_i_pregs_60 : _GEN_955; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_957 = 7'h3d == io_i_rename_table_7 ? io_i_pregs_61 : _GEN_956; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_958 = 7'h3e == io_i_rename_table_7 ? io_i_pregs_62 : _GEN_957; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_959 = 7'h3f == io_i_rename_table_7 ? io_i_pregs_63 : _GEN_958; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_960 = 7'h40 == io_i_rename_table_7 ? io_i_pregs_64 : _GEN_959; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_961 = 7'h41 == io_i_rename_table_7 ? io_i_pregs_65 : _GEN_960; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_962 = 7'h42 == io_i_rename_table_7 ? io_i_pregs_66 : _GEN_961; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_963 = 7'h43 == io_i_rename_table_7 ? io_i_pregs_67 : _GEN_962; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_964 = 7'h44 == io_i_rename_table_7 ? io_i_pregs_68 : _GEN_963; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_965 = 7'h45 == io_i_rename_table_7 ? io_i_pregs_69 : _GEN_964; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_966 = 7'h46 == io_i_rename_table_7 ? io_i_pregs_70 : _GEN_965; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_967 = 7'h47 == io_i_rename_table_7 ? io_i_pregs_71 : _GEN_966; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_968 = 7'h48 == io_i_rename_table_7 ? io_i_pregs_72 : _GEN_967; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_969 = 7'h49 == io_i_rename_table_7 ? io_i_pregs_73 : _GEN_968; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_970 = 7'h4a == io_i_rename_table_7 ? io_i_pregs_74 : _GEN_969; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_971 = 7'h4b == io_i_rename_table_7 ? io_i_pregs_75 : _GEN_970; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_972 = 7'h4c == io_i_rename_table_7 ? io_i_pregs_76 : _GEN_971; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_973 = 7'h4d == io_i_rename_table_7 ? io_i_pregs_77 : _GEN_972; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_974 = 7'h4e == io_i_rename_table_7 ? io_i_pregs_78 : _GEN_973; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_975 = 7'h4f == io_i_rename_table_7 ? io_i_pregs_79 : _GEN_974; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_976 = 7'h50 == io_i_rename_table_7 ? io_i_pregs_80 : _GEN_975; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_977 = 7'h51 == io_i_rename_table_7 ? io_i_pregs_81 : _GEN_976; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_978 = 7'h52 == io_i_rename_table_7 ? io_i_pregs_82 : _GEN_977; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_979 = 7'h53 == io_i_rename_table_7 ? io_i_pregs_83 : _GEN_978; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_980 = 7'h54 == io_i_rename_table_7 ? io_i_pregs_84 : _GEN_979; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_981 = 7'h55 == io_i_rename_table_7 ? io_i_pregs_85 : _GEN_980; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_982 = 7'h56 == io_i_rename_table_7 ? io_i_pregs_86 : _GEN_981; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_983 = 7'h57 == io_i_rename_table_7 ? io_i_pregs_87 : _GEN_982; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_984 = 7'h58 == io_i_rename_table_7 ? io_i_pregs_88 : _GEN_983; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_985 = 7'h59 == io_i_rename_table_7 ? io_i_pregs_89 : _GEN_984; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_986 = 7'h5a == io_i_rename_table_7 ? io_i_pregs_90 : _GEN_985; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_987 = 7'h5b == io_i_rename_table_7 ? io_i_pregs_91 : _GEN_986; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_988 = 7'h5c == io_i_rename_table_7 ? io_i_pregs_92 : _GEN_987; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_989 = 7'h5d == io_i_rename_table_7 ? io_i_pregs_93 : _GEN_988; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_990 = 7'h5e == io_i_rename_table_7 ? io_i_pregs_94 : _GEN_989; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_991 = 7'h5f == io_i_rename_table_7 ? io_i_pregs_95 : _GEN_990; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_992 = 7'h60 == io_i_rename_table_7 ? io_i_pregs_96 : _GEN_991; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_993 = 7'h61 == io_i_rename_table_7 ? io_i_pregs_97 : _GEN_992; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_994 = 7'h62 == io_i_rename_table_7 ? io_i_pregs_98 : _GEN_993; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_995 = 7'h63 == io_i_rename_table_7 ? io_i_pregs_99 : _GEN_994; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_996 = 7'h64 == io_i_rename_table_7 ? io_i_pregs_100 : _GEN_995; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_997 = 7'h65 == io_i_rename_table_7 ? io_i_pregs_101 : _GEN_996; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_998 = 7'h66 == io_i_rename_table_7 ? io_i_pregs_102 : _GEN_997; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_999 = 7'h67 == io_i_rename_table_7 ? io_i_pregs_103 : _GEN_998; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1000 = 7'h68 == io_i_rename_table_7 ? io_i_pregs_104 : _GEN_999; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1001 = 7'h69 == io_i_rename_table_7 ? io_i_pregs_105 : _GEN_1000; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1002 = 7'h6a == io_i_rename_table_7 ? io_i_pregs_106 : _GEN_1001; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1003 = 7'h6b == io_i_rename_table_7 ? io_i_pregs_107 : _GEN_1002; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1004 = 7'h6c == io_i_rename_table_7 ? io_i_pregs_108 : _GEN_1003; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1005 = 7'h6d == io_i_rename_table_7 ? io_i_pregs_109 : _GEN_1004; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1006 = 7'h6e == io_i_rename_table_7 ? io_i_pregs_110 : _GEN_1005; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1007 = 7'h6f == io_i_rename_table_7 ? io_i_pregs_111 : _GEN_1006; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1008 = 7'h70 == io_i_rename_table_7 ? io_i_pregs_112 : _GEN_1007; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1009 = 7'h71 == io_i_rename_table_7 ? io_i_pregs_113 : _GEN_1008; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1010 = 7'h72 == io_i_rename_table_7 ? io_i_pregs_114 : _GEN_1009; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1011 = 7'h73 == io_i_rename_table_7 ? io_i_pregs_115 : _GEN_1010; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1012 = 7'h74 == io_i_rename_table_7 ? io_i_pregs_116 : _GEN_1011; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1013 = 7'h75 == io_i_rename_table_7 ? io_i_pregs_117 : _GEN_1012; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1014 = 7'h76 == io_i_rename_table_7 ? io_i_pregs_118 : _GEN_1013; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1015 = 7'h77 == io_i_rename_table_7 ? io_i_pregs_119 : _GEN_1014; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1016 = 7'h78 == io_i_rename_table_7 ? io_i_pregs_120 : _GEN_1015; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1017 = 7'h79 == io_i_rename_table_7 ? io_i_pregs_121 : _GEN_1016; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1018 = 7'h7a == io_i_rename_table_7 ? io_i_pregs_122 : _GEN_1017; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1019 = 7'h7b == io_i_rename_table_7 ? io_i_pregs_123 : _GEN_1018; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1020 = 7'h7c == io_i_rename_table_7 ? io_i_pregs_124 : _GEN_1019; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1021 = 7'h7d == io_i_rename_table_7 ? io_i_pregs_125 : _GEN_1020; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1022 = 7'h7e == io_i_rename_table_7 ? io_i_pregs_126 : _GEN_1021; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1025 = 7'h1 == io_i_rename_table_8 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1026 = 7'h2 == io_i_rename_table_8 ? io_i_pregs_2 : _GEN_1025; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1027 = 7'h3 == io_i_rename_table_8 ? io_i_pregs_3 : _GEN_1026; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1028 = 7'h4 == io_i_rename_table_8 ? io_i_pregs_4 : _GEN_1027; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1029 = 7'h5 == io_i_rename_table_8 ? io_i_pregs_5 : _GEN_1028; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1030 = 7'h6 == io_i_rename_table_8 ? io_i_pregs_6 : _GEN_1029; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1031 = 7'h7 == io_i_rename_table_8 ? io_i_pregs_7 : _GEN_1030; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1032 = 7'h8 == io_i_rename_table_8 ? io_i_pregs_8 : _GEN_1031; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1033 = 7'h9 == io_i_rename_table_8 ? io_i_pregs_9 : _GEN_1032; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1034 = 7'ha == io_i_rename_table_8 ? io_i_pregs_10 : _GEN_1033; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1035 = 7'hb == io_i_rename_table_8 ? io_i_pregs_11 : _GEN_1034; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1036 = 7'hc == io_i_rename_table_8 ? io_i_pregs_12 : _GEN_1035; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1037 = 7'hd == io_i_rename_table_8 ? io_i_pregs_13 : _GEN_1036; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1038 = 7'he == io_i_rename_table_8 ? io_i_pregs_14 : _GEN_1037; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1039 = 7'hf == io_i_rename_table_8 ? io_i_pregs_15 : _GEN_1038; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1040 = 7'h10 == io_i_rename_table_8 ? io_i_pregs_16 : _GEN_1039; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1041 = 7'h11 == io_i_rename_table_8 ? io_i_pregs_17 : _GEN_1040; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1042 = 7'h12 == io_i_rename_table_8 ? io_i_pregs_18 : _GEN_1041; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1043 = 7'h13 == io_i_rename_table_8 ? io_i_pregs_19 : _GEN_1042; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1044 = 7'h14 == io_i_rename_table_8 ? io_i_pregs_20 : _GEN_1043; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1045 = 7'h15 == io_i_rename_table_8 ? io_i_pregs_21 : _GEN_1044; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1046 = 7'h16 == io_i_rename_table_8 ? io_i_pregs_22 : _GEN_1045; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1047 = 7'h17 == io_i_rename_table_8 ? io_i_pregs_23 : _GEN_1046; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1048 = 7'h18 == io_i_rename_table_8 ? io_i_pregs_24 : _GEN_1047; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1049 = 7'h19 == io_i_rename_table_8 ? io_i_pregs_25 : _GEN_1048; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1050 = 7'h1a == io_i_rename_table_8 ? io_i_pregs_26 : _GEN_1049; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1051 = 7'h1b == io_i_rename_table_8 ? io_i_pregs_27 : _GEN_1050; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1052 = 7'h1c == io_i_rename_table_8 ? io_i_pregs_28 : _GEN_1051; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1053 = 7'h1d == io_i_rename_table_8 ? io_i_pregs_29 : _GEN_1052; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1054 = 7'h1e == io_i_rename_table_8 ? io_i_pregs_30 : _GEN_1053; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1055 = 7'h1f == io_i_rename_table_8 ? io_i_pregs_31 : _GEN_1054; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1056 = 7'h20 == io_i_rename_table_8 ? io_i_pregs_32 : _GEN_1055; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1057 = 7'h21 == io_i_rename_table_8 ? io_i_pregs_33 : _GEN_1056; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1058 = 7'h22 == io_i_rename_table_8 ? io_i_pregs_34 : _GEN_1057; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1059 = 7'h23 == io_i_rename_table_8 ? io_i_pregs_35 : _GEN_1058; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1060 = 7'h24 == io_i_rename_table_8 ? io_i_pregs_36 : _GEN_1059; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1061 = 7'h25 == io_i_rename_table_8 ? io_i_pregs_37 : _GEN_1060; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1062 = 7'h26 == io_i_rename_table_8 ? io_i_pregs_38 : _GEN_1061; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1063 = 7'h27 == io_i_rename_table_8 ? io_i_pregs_39 : _GEN_1062; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1064 = 7'h28 == io_i_rename_table_8 ? io_i_pregs_40 : _GEN_1063; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1065 = 7'h29 == io_i_rename_table_8 ? io_i_pregs_41 : _GEN_1064; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1066 = 7'h2a == io_i_rename_table_8 ? io_i_pregs_42 : _GEN_1065; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1067 = 7'h2b == io_i_rename_table_8 ? io_i_pregs_43 : _GEN_1066; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1068 = 7'h2c == io_i_rename_table_8 ? io_i_pregs_44 : _GEN_1067; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1069 = 7'h2d == io_i_rename_table_8 ? io_i_pregs_45 : _GEN_1068; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1070 = 7'h2e == io_i_rename_table_8 ? io_i_pregs_46 : _GEN_1069; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1071 = 7'h2f == io_i_rename_table_8 ? io_i_pregs_47 : _GEN_1070; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1072 = 7'h30 == io_i_rename_table_8 ? io_i_pregs_48 : _GEN_1071; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1073 = 7'h31 == io_i_rename_table_8 ? io_i_pregs_49 : _GEN_1072; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1074 = 7'h32 == io_i_rename_table_8 ? io_i_pregs_50 : _GEN_1073; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1075 = 7'h33 == io_i_rename_table_8 ? io_i_pregs_51 : _GEN_1074; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1076 = 7'h34 == io_i_rename_table_8 ? io_i_pregs_52 : _GEN_1075; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1077 = 7'h35 == io_i_rename_table_8 ? io_i_pregs_53 : _GEN_1076; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1078 = 7'h36 == io_i_rename_table_8 ? io_i_pregs_54 : _GEN_1077; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1079 = 7'h37 == io_i_rename_table_8 ? io_i_pregs_55 : _GEN_1078; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1080 = 7'h38 == io_i_rename_table_8 ? io_i_pregs_56 : _GEN_1079; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1081 = 7'h39 == io_i_rename_table_8 ? io_i_pregs_57 : _GEN_1080; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1082 = 7'h3a == io_i_rename_table_8 ? io_i_pregs_58 : _GEN_1081; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1083 = 7'h3b == io_i_rename_table_8 ? io_i_pregs_59 : _GEN_1082; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1084 = 7'h3c == io_i_rename_table_8 ? io_i_pregs_60 : _GEN_1083; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1085 = 7'h3d == io_i_rename_table_8 ? io_i_pregs_61 : _GEN_1084; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1086 = 7'h3e == io_i_rename_table_8 ? io_i_pregs_62 : _GEN_1085; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1087 = 7'h3f == io_i_rename_table_8 ? io_i_pregs_63 : _GEN_1086; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1088 = 7'h40 == io_i_rename_table_8 ? io_i_pregs_64 : _GEN_1087; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1089 = 7'h41 == io_i_rename_table_8 ? io_i_pregs_65 : _GEN_1088; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1090 = 7'h42 == io_i_rename_table_8 ? io_i_pregs_66 : _GEN_1089; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1091 = 7'h43 == io_i_rename_table_8 ? io_i_pregs_67 : _GEN_1090; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1092 = 7'h44 == io_i_rename_table_8 ? io_i_pregs_68 : _GEN_1091; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1093 = 7'h45 == io_i_rename_table_8 ? io_i_pregs_69 : _GEN_1092; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1094 = 7'h46 == io_i_rename_table_8 ? io_i_pregs_70 : _GEN_1093; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1095 = 7'h47 == io_i_rename_table_8 ? io_i_pregs_71 : _GEN_1094; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1096 = 7'h48 == io_i_rename_table_8 ? io_i_pregs_72 : _GEN_1095; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1097 = 7'h49 == io_i_rename_table_8 ? io_i_pregs_73 : _GEN_1096; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1098 = 7'h4a == io_i_rename_table_8 ? io_i_pregs_74 : _GEN_1097; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1099 = 7'h4b == io_i_rename_table_8 ? io_i_pregs_75 : _GEN_1098; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1100 = 7'h4c == io_i_rename_table_8 ? io_i_pregs_76 : _GEN_1099; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1101 = 7'h4d == io_i_rename_table_8 ? io_i_pregs_77 : _GEN_1100; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1102 = 7'h4e == io_i_rename_table_8 ? io_i_pregs_78 : _GEN_1101; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1103 = 7'h4f == io_i_rename_table_8 ? io_i_pregs_79 : _GEN_1102; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1104 = 7'h50 == io_i_rename_table_8 ? io_i_pregs_80 : _GEN_1103; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1105 = 7'h51 == io_i_rename_table_8 ? io_i_pregs_81 : _GEN_1104; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1106 = 7'h52 == io_i_rename_table_8 ? io_i_pregs_82 : _GEN_1105; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1107 = 7'h53 == io_i_rename_table_8 ? io_i_pregs_83 : _GEN_1106; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1108 = 7'h54 == io_i_rename_table_8 ? io_i_pregs_84 : _GEN_1107; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1109 = 7'h55 == io_i_rename_table_8 ? io_i_pregs_85 : _GEN_1108; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1110 = 7'h56 == io_i_rename_table_8 ? io_i_pregs_86 : _GEN_1109; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1111 = 7'h57 == io_i_rename_table_8 ? io_i_pregs_87 : _GEN_1110; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1112 = 7'h58 == io_i_rename_table_8 ? io_i_pregs_88 : _GEN_1111; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1113 = 7'h59 == io_i_rename_table_8 ? io_i_pregs_89 : _GEN_1112; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1114 = 7'h5a == io_i_rename_table_8 ? io_i_pregs_90 : _GEN_1113; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1115 = 7'h5b == io_i_rename_table_8 ? io_i_pregs_91 : _GEN_1114; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1116 = 7'h5c == io_i_rename_table_8 ? io_i_pregs_92 : _GEN_1115; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1117 = 7'h5d == io_i_rename_table_8 ? io_i_pregs_93 : _GEN_1116; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1118 = 7'h5e == io_i_rename_table_8 ? io_i_pregs_94 : _GEN_1117; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1119 = 7'h5f == io_i_rename_table_8 ? io_i_pregs_95 : _GEN_1118; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1120 = 7'h60 == io_i_rename_table_8 ? io_i_pregs_96 : _GEN_1119; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1121 = 7'h61 == io_i_rename_table_8 ? io_i_pregs_97 : _GEN_1120; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1122 = 7'h62 == io_i_rename_table_8 ? io_i_pregs_98 : _GEN_1121; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1123 = 7'h63 == io_i_rename_table_8 ? io_i_pregs_99 : _GEN_1122; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1124 = 7'h64 == io_i_rename_table_8 ? io_i_pregs_100 : _GEN_1123; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1125 = 7'h65 == io_i_rename_table_8 ? io_i_pregs_101 : _GEN_1124; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1126 = 7'h66 == io_i_rename_table_8 ? io_i_pregs_102 : _GEN_1125; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1127 = 7'h67 == io_i_rename_table_8 ? io_i_pregs_103 : _GEN_1126; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1128 = 7'h68 == io_i_rename_table_8 ? io_i_pregs_104 : _GEN_1127; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1129 = 7'h69 == io_i_rename_table_8 ? io_i_pregs_105 : _GEN_1128; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1130 = 7'h6a == io_i_rename_table_8 ? io_i_pregs_106 : _GEN_1129; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1131 = 7'h6b == io_i_rename_table_8 ? io_i_pregs_107 : _GEN_1130; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1132 = 7'h6c == io_i_rename_table_8 ? io_i_pregs_108 : _GEN_1131; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1133 = 7'h6d == io_i_rename_table_8 ? io_i_pregs_109 : _GEN_1132; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1134 = 7'h6e == io_i_rename_table_8 ? io_i_pregs_110 : _GEN_1133; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1135 = 7'h6f == io_i_rename_table_8 ? io_i_pregs_111 : _GEN_1134; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1136 = 7'h70 == io_i_rename_table_8 ? io_i_pregs_112 : _GEN_1135; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1137 = 7'h71 == io_i_rename_table_8 ? io_i_pregs_113 : _GEN_1136; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1138 = 7'h72 == io_i_rename_table_8 ? io_i_pregs_114 : _GEN_1137; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1139 = 7'h73 == io_i_rename_table_8 ? io_i_pregs_115 : _GEN_1138; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1140 = 7'h74 == io_i_rename_table_8 ? io_i_pregs_116 : _GEN_1139; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1141 = 7'h75 == io_i_rename_table_8 ? io_i_pregs_117 : _GEN_1140; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1142 = 7'h76 == io_i_rename_table_8 ? io_i_pregs_118 : _GEN_1141; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1143 = 7'h77 == io_i_rename_table_8 ? io_i_pregs_119 : _GEN_1142; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1144 = 7'h78 == io_i_rename_table_8 ? io_i_pregs_120 : _GEN_1143; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1145 = 7'h79 == io_i_rename_table_8 ? io_i_pregs_121 : _GEN_1144; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1146 = 7'h7a == io_i_rename_table_8 ? io_i_pregs_122 : _GEN_1145; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1147 = 7'h7b == io_i_rename_table_8 ? io_i_pregs_123 : _GEN_1146; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1148 = 7'h7c == io_i_rename_table_8 ? io_i_pregs_124 : _GEN_1147; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1149 = 7'h7d == io_i_rename_table_8 ? io_i_pregs_125 : _GEN_1148; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1150 = 7'h7e == io_i_rename_table_8 ? io_i_pregs_126 : _GEN_1149; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1153 = 7'h1 == io_i_rename_table_9 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1154 = 7'h2 == io_i_rename_table_9 ? io_i_pregs_2 : _GEN_1153; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1155 = 7'h3 == io_i_rename_table_9 ? io_i_pregs_3 : _GEN_1154; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1156 = 7'h4 == io_i_rename_table_9 ? io_i_pregs_4 : _GEN_1155; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1157 = 7'h5 == io_i_rename_table_9 ? io_i_pregs_5 : _GEN_1156; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1158 = 7'h6 == io_i_rename_table_9 ? io_i_pregs_6 : _GEN_1157; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1159 = 7'h7 == io_i_rename_table_9 ? io_i_pregs_7 : _GEN_1158; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1160 = 7'h8 == io_i_rename_table_9 ? io_i_pregs_8 : _GEN_1159; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1161 = 7'h9 == io_i_rename_table_9 ? io_i_pregs_9 : _GEN_1160; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1162 = 7'ha == io_i_rename_table_9 ? io_i_pregs_10 : _GEN_1161; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1163 = 7'hb == io_i_rename_table_9 ? io_i_pregs_11 : _GEN_1162; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1164 = 7'hc == io_i_rename_table_9 ? io_i_pregs_12 : _GEN_1163; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1165 = 7'hd == io_i_rename_table_9 ? io_i_pregs_13 : _GEN_1164; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1166 = 7'he == io_i_rename_table_9 ? io_i_pregs_14 : _GEN_1165; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1167 = 7'hf == io_i_rename_table_9 ? io_i_pregs_15 : _GEN_1166; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1168 = 7'h10 == io_i_rename_table_9 ? io_i_pregs_16 : _GEN_1167; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1169 = 7'h11 == io_i_rename_table_9 ? io_i_pregs_17 : _GEN_1168; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1170 = 7'h12 == io_i_rename_table_9 ? io_i_pregs_18 : _GEN_1169; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1171 = 7'h13 == io_i_rename_table_9 ? io_i_pregs_19 : _GEN_1170; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1172 = 7'h14 == io_i_rename_table_9 ? io_i_pregs_20 : _GEN_1171; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1173 = 7'h15 == io_i_rename_table_9 ? io_i_pregs_21 : _GEN_1172; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1174 = 7'h16 == io_i_rename_table_9 ? io_i_pregs_22 : _GEN_1173; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1175 = 7'h17 == io_i_rename_table_9 ? io_i_pregs_23 : _GEN_1174; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1176 = 7'h18 == io_i_rename_table_9 ? io_i_pregs_24 : _GEN_1175; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1177 = 7'h19 == io_i_rename_table_9 ? io_i_pregs_25 : _GEN_1176; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1178 = 7'h1a == io_i_rename_table_9 ? io_i_pregs_26 : _GEN_1177; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1179 = 7'h1b == io_i_rename_table_9 ? io_i_pregs_27 : _GEN_1178; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1180 = 7'h1c == io_i_rename_table_9 ? io_i_pregs_28 : _GEN_1179; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1181 = 7'h1d == io_i_rename_table_9 ? io_i_pregs_29 : _GEN_1180; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1182 = 7'h1e == io_i_rename_table_9 ? io_i_pregs_30 : _GEN_1181; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1183 = 7'h1f == io_i_rename_table_9 ? io_i_pregs_31 : _GEN_1182; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1184 = 7'h20 == io_i_rename_table_9 ? io_i_pregs_32 : _GEN_1183; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1185 = 7'h21 == io_i_rename_table_9 ? io_i_pregs_33 : _GEN_1184; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1186 = 7'h22 == io_i_rename_table_9 ? io_i_pregs_34 : _GEN_1185; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1187 = 7'h23 == io_i_rename_table_9 ? io_i_pregs_35 : _GEN_1186; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1188 = 7'h24 == io_i_rename_table_9 ? io_i_pregs_36 : _GEN_1187; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1189 = 7'h25 == io_i_rename_table_9 ? io_i_pregs_37 : _GEN_1188; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1190 = 7'h26 == io_i_rename_table_9 ? io_i_pregs_38 : _GEN_1189; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1191 = 7'h27 == io_i_rename_table_9 ? io_i_pregs_39 : _GEN_1190; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1192 = 7'h28 == io_i_rename_table_9 ? io_i_pregs_40 : _GEN_1191; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1193 = 7'h29 == io_i_rename_table_9 ? io_i_pregs_41 : _GEN_1192; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1194 = 7'h2a == io_i_rename_table_9 ? io_i_pregs_42 : _GEN_1193; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1195 = 7'h2b == io_i_rename_table_9 ? io_i_pregs_43 : _GEN_1194; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1196 = 7'h2c == io_i_rename_table_9 ? io_i_pregs_44 : _GEN_1195; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1197 = 7'h2d == io_i_rename_table_9 ? io_i_pregs_45 : _GEN_1196; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1198 = 7'h2e == io_i_rename_table_9 ? io_i_pregs_46 : _GEN_1197; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1199 = 7'h2f == io_i_rename_table_9 ? io_i_pregs_47 : _GEN_1198; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1200 = 7'h30 == io_i_rename_table_9 ? io_i_pregs_48 : _GEN_1199; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1201 = 7'h31 == io_i_rename_table_9 ? io_i_pregs_49 : _GEN_1200; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1202 = 7'h32 == io_i_rename_table_9 ? io_i_pregs_50 : _GEN_1201; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1203 = 7'h33 == io_i_rename_table_9 ? io_i_pregs_51 : _GEN_1202; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1204 = 7'h34 == io_i_rename_table_9 ? io_i_pregs_52 : _GEN_1203; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1205 = 7'h35 == io_i_rename_table_9 ? io_i_pregs_53 : _GEN_1204; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1206 = 7'h36 == io_i_rename_table_9 ? io_i_pregs_54 : _GEN_1205; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1207 = 7'h37 == io_i_rename_table_9 ? io_i_pregs_55 : _GEN_1206; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1208 = 7'h38 == io_i_rename_table_9 ? io_i_pregs_56 : _GEN_1207; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1209 = 7'h39 == io_i_rename_table_9 ? io_i_pregs_57 : _GEN_1208; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1210 = 7'h3a == io_i_rename_table_9 ? io_i_pregs_58 : _GEN_1209; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1211 = 7'h3b == io_i_rename_table_9 ? io_i_pregs_59 : _GEN_1210; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1212 = 7'h3c == io_i_rename_table_9 ? io_i_pregs_60 : _GEN_1211; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1213 = 7'h3d == io_i_rename_table_9 ? io_i_pregs_61 : _GEN_1212; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1214 = 7'h3e == io_i_rename_table_9 ? io_i_pregs_62 : _GEN_1213; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1215 = 7'h3f == io_i_rename_table_9 ? io_i_pregs_63 : _GEN_1214; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1216 = 7'h40 == io_i_rename_table_9 ? io_i_pregs_64 : _GEN_1215; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1217 = 7'h41 == io_i_rename_table_9 ? io_i_pregs_65 : _GEN_1216; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1218 = 7'h42 == io_i_rename_table_9 ? io_i_pregs_66 : _GEN_1217; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1219 = 7'h43 == io_i_rename_table_9 ? io_i_pregs_67 : _GEN_1218; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1220 = 7'h44 == io_i_rename_table_9 ? io_i_pregs_68 : _GEN_1219; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1221 = 7'h45 == io_i_rename_table_9 ? io_i_pregs_69 : _GEN_1220; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1222 = 7'h46 == io_i_rename_table_9 ? io_i_pregs_70 : _GEN_1221; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1223 = 7'h47 == io_i_rename_table_9 ? io_i_pregs_71 : _GEN_1222; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1224 = 7'h48 == io_i_rename_table_9 ? io_i_pregs_72 : _GEN_1223; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1225 = 7'h49 == io_i_rename_table_9 ? io_i_pregs_73 : _GEN_1224; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1226 = 7'h4a == io_i_rename_table_9 ? io_i_pregs_74 : _GEN_1225; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1227 = 7'h4b == io_i_rename_table_9 ? io_i_pregs_75 : _GEN_1226; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1228 = 7'h4c == io_i_rename_table_9 ? io_i_pregs_76 : _GEN_1227; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1229 = 7'h4d == io_i_rename_table_9 ? io_i_pregs_77 : _GEN_1228; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1230 = 7'h4e == io_i_rename_table_9 ? io_i_pregs_78 : _GEN_1229; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1231 = 7'h4f == io_i_rename_table_9 ? io_i_pregs_79 : _GEN_1230; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1232 = 7'h50 == io_i_rename_table_9 ? io_i_pregs_80 : _GEN_1231; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1233 = 7'h51 == io_i_rename_table_9 ? io_i_pregs_81 : _GEN_1232; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1234 = 7'h52 == io_i_rename_table_9 ? io_i_pregs_82 : _GEN_1233; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1235 = 7'h53 == io_i_rename_table_9 ? io_i_pregs_83 : _GEN_1234; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1236 = 7'h54 == io_i_rename_table_9 ? io_i_pregs_84 : _GEN_1235; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1237 = 7'h55 == io_i_rename_table_9 ? io_i_pregs_85 : _GEN_1236; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1238 = 7'h56 == io_i_rename_table_9 ? io_i_pregs_86 : _GEN_1237; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1239 = 7'h57 == io_i_rename_table_9 ? io_i_pregs_87 : _GEN_1238; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1240 = 7'h58 == io_i_rename_table_9 ? io_i_pregs_88 : _GEN_1239; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1241 = 7'h59 == io_i_rename_table_9 ? io_i_pregs_89 : _GEN_1240; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1242 = 7'h5a == io_i_rename_table_9 ? io_i_pregs_90 : _GEN_1241; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1243 = 7'h5b == io_i_rename_table_9 ? io_i_pregs_91 : _GEN_1242; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1244 = 7'h5c == io_i_rename_table_9 ? io_i_pregs_92 : _GEN_1243; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1245 = 7'h5d == io_i_rename_table_9 ? io_i_pregs_93 : _GEN_1244; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1246 = 7'h5e == io_i_rename_table_9 ? io_i_pregs_94 : _GEN_1245; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1247 = 7'h5f == io_i_rename_table_9 ? io_i_pregs_95 : _GEN_1246; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1248 = 7'h60 == io_i_rename_table_9 ? io_i_pregs_96 : _GEN_1247; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1249 = 7'h61 == io_i_rename_table_9 ? io_i_pregs_97 : _GEN_1248; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1250 = 7'h62 == io_i_rename_table_9 ? io_i_pregs_98 : _GEN_1249; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1251 = 7'h63 == io_i_rename_table_9 ? io_i_pregs_99 : _GEN_1250; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1252 = 7'h64 == io_i_rename_table_9 ? io_i_pregs_100 : _GEN_1251; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1253 = 7'h65 == io_i_rename_table_9 ? io_i_pregs_101 : _GEN_1252; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1254 = 7'h66 == io_i_rename_table_9 ? io_i_pregs_102 : _GEN_1253; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1255 = 7'h67 == io_i_rename_table_9 ? io_i_pregs_103 : _GEN_1254; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1256 = 7'h68 == io_i_rename_table_9 ? io_i_pregs_104 : _GEN_1255; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1257 = 7'h69 == io_i_rename_table_9 ? io_i_pregs_105 : _GEN_1256; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1258 = 7'h6a == io_i_rename_table_9 ? io_i_pregs_106 : _GEN_1257; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1259 = 7'h6b == io_i_rename_table_9 ? io_i_pregs_107 : _GEN_1258; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1260 = 7'h6c == io_i_rename_table_9 ? io_i_pregs_108 : _GEN_1259; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1261 = 7'h6d == io_i_rename_table_9 ? io_i_pregs_109 : _GEN_1260; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1262 = 7'h6e == io_i_rename_table_9 ? io_i_pregs_110 : _GEN_1261; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1263 = 7'h6f == io_i_rename_table_9 ? io_i_pregs_111 : _GEN_1262; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1264 = 7'h70 == io_i_rename_table_9 ? io_i_pregs_112 : _GEN_1263; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1265 = 7'h71 == io_i_rename_table_9 ? io_i_pregs_113 : _GEN_1264; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1266 = 7'h72 == io_i_rename_table_9 ? io_i_pregs_114 : _GEN_1265; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1267 = 7'h73 == io_i_rename_table_9 ? io_i_pregs_115 : _GEN_1266; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1268 = 7'h74 == io_i_rename_table_9 ? io_i_pregs_116 : _GEN_1267; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1269 = 7'h75 == io_i_rename_table_9 ? io_i_pregs_117 : _GEN_1268; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1270 = 7'h76 == io_i_rename_table_9 ? io_i_pregs_118 : _GEN_1269; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1271 = 7'h77 == io_i_rename_table_9 ? io_i_pregs_119 : _GEN_1270; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1272 = 7'h78 == io_i_rename_table_9 ? io_i_pregs_120 : _GEN_1271; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1273 = 7'h79 == io_i_rename_table_9 ? io_i_pregs_121 : _GEN_1272; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1274 = 7'h7a == io_i_rename_table_9 ? io_i_pregs_122 : _GEN_1273; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1275 = 7'h7b == io_i_rename_table_9 ? io_i_pregs_123 : _GEN_1274; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1276 = 7'h7c == io_i_rename_table_9 ? io_i_pregs_124 : _GEN_1275; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1277 = 7'h7d == io_i_rename_table_9 ? io_i_pregs_125 : _GEN_1276; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1278 = 7'h7e == io_i_rename_table_9 ? io_i_pregs_126 : _GEN_1277; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1281 = 7'h1 == io_i_rename_table_10 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1282 = 7'h2 == io_i_rename_table_10 ? io_i_pregs_2 : _GEN_1281; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1283 = 7'h3 == io_i_rename_table_10 ? io_i_pregs_3 : _GEN_1282; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1284 = 7'h4 == io_i_rename_table_10 ? io_i_pregs_4 : _GEN_1283; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1285 = 7'h5 == io_i_rename_table_10 ? io_i_pregs_5 : _GEN_1284; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1286 = 7'h6 == io_i_rename_table_10 ? io_i_pregs_6 : _GEN_1285; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1287 = 7'h7 == io_i_rename_table_10 ? io_i_pregs_7 : _GEN_1286; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1288 = 7'h8 == io_i_rename_table_10 ? io_i_pregs_8 : _GEN_1287; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1289 = 7'h9 == io_i_rename_table_10 ? io_i_pregs_9 : _GEN_1288; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1290 = 7'ha == io_i_rename_table_10 ? io_i_pregs_10 : _GEN_1289; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1291 = 7'hb == io_i_rename_table_10 ? io_i_pregs_11 : _GEN_1290; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1292 = 7'hc == io_i_rename_table_10 ? io_i_pregs_12 : _GEN_1291; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1293 = 7'hd == io_i_rename_table_10 ? io_i_pregs_13 : _GEN_1292; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1294 = 7'he == io_i_rename_table_10 ? io_i_pregs_14 : _GEN_1293; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1295 = 7'hf == io_i_rename_table_10 ? io_i_pregs_15 : _GEN_1294; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1296 = 7'h10 == io_i_rename_table_10 ? io_i_pregs_16 : _GEN_1295; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1297 = 7'h11 == io_i_rename_table_10 ? io_i_pregs_17 : _GEN_1296; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1298 = 7'h12 == io_i_rename_table_10 ? io_i_pregs_18 : _GEN_1297; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1299 = 7'h13 == io_i_rename_table_10 ? io_i_pregs_19 : _GEN_1298; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1300 = 7'h14 == io_i_rename_table_10 ? io_i_pregs_20 : _GEN_1299; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1301 = 7'h15 == io_i_rename_table_10 ? io_i_pregs_21 : _GEN_1300; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1302 = 7'h16 == io_i_rename_table_10 ? io_i_pregs_22 : _GEN_1301; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1303 = 7'h17 == io_i_rename_table_10 ? io_i_pregs_23 : _GEN_1302; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1304 = 7'h18 == io_i_rename_table_10 ? io_i_pregs_24 : _GEN_1303; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1305 = 7'h19 == io_i_rename_table_10 ? io_i_pregs_25 : _GEN_1304; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1306 = 7'h1a == io_i_rename_table_10 ? io_i_pregs_26 : _GEN_1305; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1307 = 7'h1b == io_i_rename_table_10 ? io_i_pregs_27 : _GEN_1306; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1308 = 7'h1c == io_i_rename_table_10 ? io_i_pregs_28 : _GEN_1307; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1309 = 7'h1d == io_i_rename_table_10 ? io_i_pregs_29 : _GEN_1308; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1310 = 7'h1e == io_i_rename_table_10 ? io_i_pregs_30 : _GEN_1309; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1311 = 7'h1f == io_i_rename_table_10 ? io_i_pregs_31 : _GEN_1310; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1312 = 7'h20 == io_i_rename_table_10 ? io_i_pregs_32 : _GEN_1311; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1313 = 7'h21 == io_i_rename_table_10 ? io_i_pregs_33 : _GEN_1312; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1314 = 7'h22 == io_i_rename_table_10 ? io_i_pregs_34 : _GEN_1313; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1315 = 7'h23 == io_i_rename_table_10 ? io_i_pregs_35 : _GEN_1314; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1316 = 7'h24 == io_i_rename_table_10 ? io_i_pregs_36 : _GEN_1315; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1317 = 7'h25 == io_i_rename_table_10 ? io_i_pregs_37 : _GEN_1316; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1318 = 7'h26 == io_i_rename_table_10 ? io_i_pregs_38 : _GEN_1317; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1319 = 7'h27 == io_i_rename_table_10 ? io_i_pregs_39 : _GEN_1318; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1320 = 7'h28 == io_i_rename_table_10 ? io_i_pregs_40 : _GEN_1319; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1321 = 7'h29 == io_i_rename_table_10 ? io_i_pregs_41 : _GEN_1320; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1322 = 7'h2a == io_i_rename_table_10 ? io_i_pregs_42 : _GEN_1321; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1323 = 7'h2b == io_i_rename_table_10 ? io_i_pregs_43 : _GEN_1322; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1324 = 7'h2c == io_i_rename_table_10 ? io_i_pregs_44 : _GEN_1323; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1325 = 7'h2d == io_i_rename_table_10 ? io_i_pregs_45 : _GEN_1324; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1326 = 7'h2e == io_i_rename_table_10 ? io_i_pregs_46 : _GEN_1325; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1327 = 7'h2f == io_i_rename_table_10 ? io_i_pregs_47 : _GEN_1326; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1328 = 7'h30 == io_i_rename_table_10 ? io_i_pregs_48 : _GEN_1327; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1329 = 7'h31 == io_i_rename_table_10 ? io_i_pregs_49 : _GEN_1328; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1330 = 7'h32 == io_i_rename_table_10 ? io_i_pregs_50 : _GEN_1329; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1331 = 7'h33 == io_i_rename_table_10 ? io_i_pregs_51 : _GEN_1330; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1332 = 7'h34 == io_i_rename_table_10 ? io_i_pregs_52 : _GEN_1331; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1333 = 7'h35 == io_i_rename_table_10 ? io_i_pregs_53 : _GEN_1332; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1334 = 7'h36 == io_i_rename_table_10 ? io_i_pregs_54 : _GEN_1333; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1335 = 7'h37 == io_i_rename_table_10 ? io_i_pregs_55 : _GEN_1334; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1336 = 7'h38 == io_i_rename_table_10 ? io_i_pregs_56 : _GEN_1335; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1337 = 7'h39 == io_i_rename_table_10 ? io_i_pregs_57 : _GEN_1336; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1338 = 7'h3a == io_i_rename_table_10 ? io_i_pregs_58 : _GEN_1337; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1339 = 7'h3b == io_i_rename_table_10 ? io_i_pregs_59 : _GEN_1338; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1340 = 7'h3c == io_i_rename_table_10 ? io_i_pregs_60 : _GEN_1339; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1341 = 7'h3d == io_i_rename_table_10 ? io_i_pregs_61 : _GEN_1340; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1342 = 7'h3e == io_i_rename_table_10 ? io_i_pregs_62 : _GEN_1341; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1343 = 7'h3f == io_i_rename_table_10 ? io_i_pregs_63 : _GEN_1342; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1344 = 7'h40 == io_i_rename_table_10 ? io_i_pregs_64 : _GEN_1343; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1345 = 7'h41 == io_i_rename_table_10 ? io_i_pregs_65 : _GEN_1344; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1346 = 7'h42 == io_i_rename_table_10 ? io_i_pregs_66 : _GEN_1345; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1347 = 7'h43 == io_i_rename_table_10 ? io_i_pregs_67 : _GEN_1346; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1348 = 7'h44 == io_i_rename_table_10 ? io_i_pregs_68 : _GEN_1347; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1349 = 7'h45 == io_i_rename_table_10 ? io_i_pregs_69 : _GEN_1348; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1350 = 7'h46 == io_i_rename_table_10 ? io_i_pregs_70 : _GEN_1349; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1351 = 7'h47 == io_i_rename_table_10 ? io_i_pregs_71 : _GEN_1350; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1352 = 7'h48 == io_i_rename_table_10 ? io_i_pregs_72 : _GEN_1351; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1353 = 7'h49 == io_i_rename_table_10 ? io_i_pregs_73 : _GEN_1352; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1354 = 7'h4a == io_i_rename_table_10 ? io_i_pregs_74 : _GEN_1353; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1355 = 7'h4b == io_i_rename_table_10 ? io_i_pregs_75 : _GEN_1354; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1356 = 7'h4c == io_i_rename_table_10 ? io_i_pregs_76 : _GEN_1355; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1357 = 7'h4d == io_i_rename_table_10 ? io_i_pregs_77 : _GEN_1356; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1358 = 7'h4e == io_i_rename_table_10 ? io_i_pregs_78 : _GEN_1357; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1359 = 7'h4f == io_i_rename_table_10 ? io_i_pregs_79 : _GEN_1358; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1360 = 7'h50 == io_i_rename_table_10 ? io_i_pregs_80 : _GEN_1359; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1361 = 7'h51 == io_i_rename_table_10 ? io_i_pregs_81 : _GEN_1360; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1362 = 7'h52 == io_i_rename_table_10 ? io_i_pregs_82 : _GEN_1361; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1363 = 7'h53 == io_i_rename_table_10 ? io_i_pregs_83 : _GEN_1362; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1364 = 7'h54 == io_i_rename_table_10 ? io_i_pregs_84 : _GEN_1363; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1365 = 7'h55 == io_i_rename_table_10 ? io_i_pregs_85 : _GEN_1364; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1366 = 7'h56 == io_i_rename_table_10 ? io_i_pregs_86 : _GEN_1365; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1367 = 7'h57 == io_i_rename_table_10 ? io_i_pregs_87 : _GEN_1366; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1368 = 7'h58 == io_i_rename_table_10 ? io_i_pregs_88 : _GEN_1367; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1369 = 7'h59 == io_i_rename_table_10 ? io_i_pregs_89 : _GEN_1368; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1370 = 7'h5a == io_i_rename_table_10 ? io_i_pregs_90 : _GEN_1369; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1371 = 7'h5b == io_i_rename_table_10 ? io_i_pregs_91 : _GEN_1370; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1372 = 7'h5c == io_i_rename_table_10 ? io_i_pregs_92 : _GEN_1371; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1373 = 7'h5d == io_i_rename_table_10 ? io_i_pregs_93 : _GEN_1372; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1374 = 7'h5e == io_i_rename_table_10 ? io_i_pregs_94 : _GEN_1373; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1375 = 7'h5f == io_i_rename_table_10 ? io_i_pregs_95 : _GEN_1374; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1376 = 7'h60 == io_i_rename_table_10 ? io_i_pregs_96 : _GEN_1375; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1377 = 7'h61 == io_i_rename_table_10 ? io_i_pregs_97 : _GEN_1376; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1378 = 7'h62 == io_i_rename_table_10 ? io_i_pregs_98 : _GEN_1377; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1379 = 7'h63 == io_i_rename_table_10 ? io_i_pregs_99 : _GEN_1378; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1380 = 7'h64 == io_i_rename_table_10 ? io_i_pregs_100 : _GEN_1379; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1381 = 7'h65 == io_i_rename_table_10 ? io_i_pregs_101 : _GEN_1380; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1382 = 7'h66 == io_i_rename_table_10 ? io_i_pregs_102 : _GEN_1381; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1383 = 7'h67 == io_i_rename_table_10 ? io_i_pregs_103 : _GEN_1382; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1384 = 7'h68 == io_i_rename_table_10 ? io_i_pregs_104 : _GEN_1383; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1385 = 7'h69 == io_i_rename_table_10 ? io_i_pregs_105 : _GEN_1384; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1386 = 7'h6a == io_i_rename_table_10 ? io_i_pregs_106 : _GEN_1385; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1387 = 7'h6b == io_i_rename_table_10 ? io_i_pregs_107 : _GEN_1386; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1388 = 7'h6c == io_i_rename_table_10 ? io_i_pregs_108 : _GEN_1387; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1389 = 7'h6d == io_i_rename_table_10 ? io_i_pregs_109 : _GEN_1388; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1390 = 7'h6e == io_i_rename_table_10 ? io_i_pregs_110 : _GEN_1389; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1391 = 7'h6f == io_i_rename_table_10 ? io_i_pregs_111 : _GEN_1390; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1392 = 7'h70 == io_i_rename_table_10 ? io_i_pregs_112 : _GEN_1391; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1393 = 7'h71 == io_i_rename_table_10 ? io_i_pregs_113 : _GEN_1392; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1394 = 7'h72 == io_i_rename_table_10 ? io_i_pregs_114 : _GEN_1393; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1395 = 7'h73 == io_i_rename_table_10 ? io_i_pregs_115 : _GEN_1394; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1396 = 7'h74 == io_i_rename_table_10 ? io_i_pregs_116 : _GEN_1395; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1397 = 7'h75 == io_i_rename_table_10 ? io_i_pregs_117 : _GEN_1396; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1398 = 7'h76 == io_i_rename_table_10 ? io_i_pregs_118 : _GEN_1397; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1399 = 7'h77 == io_i_rename_table_10 ? io_i_pregs_119 : _GEN_1398; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1400 = 7'h78 == io_i_rename_table_10 ? io_i_pregs_120 : _GEN_1399; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1401 = 7'h79 == io_i_rename_table_10 ? io_i_pregs_121 : _GEN_1400; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1402 = 7'h7a == io_i_rename_table_10 ? io_i_pregs_122 : _GEN_1401; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1403 = 7'h7b == io_i_rename_table_10 ? io_i_pregs_123 : _GEN_1402; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1404 = 7'h7c == io_i_rename_table_10 ? io_i_pregs_124 : _GEN_1403; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1405 = 7'h7d == io_i_rename_table_10 ? io_i_pregs_125 : _GEN_1404; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1406 = 7'h7e == io_i_rename_table_10 ? io_i_pregs_126 : _GEN_1405; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1409 = 7'h1 == io_i_rename_table_11 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1410 = 7'h2 == io_i_rename_table_11 ? io_i_pregs_2 : _GEN_1409; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1411 = 7'h3 == io_i_rename_table_11 ? io_i_pregs_3 : _GEN_1410; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1412 = 7'h4 == io_i_rename_table_11 ? io_i_pregs_4 : _GEN_1411; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1413 = 7'h5 == io_i_rename_table_11 ? io_i_pregs_5 : _GEN_1412; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1414 = 7'h6 == io_i_rename_table_11 ? io_i_pregs_6 : _GEN_1413; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1415 = 7'h7 == io_i_rename_table_11 ? io_i_pregs_7 : _GEN_1414; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1416 = 7'h8 == io_i_rename_table_11 ? io_i_pregs_8 : _GEN_1415; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1417 = 7'h9 == io_i_rename_table_11 ? io_i_pregs_9 : _GEN_1416; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1418 = 7'ha == io_i_rename_table_11 ? io_i_pregs_10 : _GEN_1417; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1419 = 7'hb == io_i_rename_table_11 ? io_i_pregs_11 : _GEN_1418; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1420 = 7'hc == io_i_rename_table_11 ? io_i_pregs_12 : _GEN_1419; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1421 = 7'hd == io_i_rename_table_11 ? io_i_pregs_13 : _GEN_1420; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1422 = 7'he == io_i_rename_table_11 ? io_i_pregs_14 : _GEN_1421; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1423 = 7'hf == io_i_rename_table_11 ? io_i_pregs_15 : _GEN_1422; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1424 = 7'h10 == io_i_rename_table_11 ? io_i_pregs_16 : _GEN_1423; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1425 = 7'h11 == io_i_rename_table_11 ? io_i_pregs_17 : _GEN_1424; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1426 = 7'h12 == io_i_rename_table_11 ? io_i_pregs_18 : _GEN_1425; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1427 = 7'h13 == io_i_rename_table_11 ? io_i_pregs_19 : _GEN_1426; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1428 = 7'h14 == io_i_rename_table_11 ? io_i_pregs_20 : _GEN_1427; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1429 = 7'h15 == io_i_rename_table_11 ? io_i_pregs_21 : _GEN_1428; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1430 = 7'h16 == io_i_rename_table_11 ? io_i_pregs_22 : _GEN_1429; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1431 = 7'h17 == io_i_rename_table_11 ? io_i_pregs_23 : _GEN_1430; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1432 = 7'h18 == io_i_rename_table_11 ? io_i_pregs_24 : _GEN_1431; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1433 = 7'h19 == io_i_rename_table_11 ? io_i_pregs_25 : _GEN_1432; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1434 = 7'h1a == io_i_rename_table_11 ? io_i_pregs_26 : _GEN_1433; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1435 = 7'h1b == io_i_rename_table_11 ? io_i_pregs_27 : _GEN_1434; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1436 = 7'h1c == io_i_rename_table_11 ? io_i_pregs_28 : _GEN_1435; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1437 = 7'h1d == io_i_rename_table_11 ? io_i_pregs_29 : _GEN_1436; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1438 = 7'h1e == io_i_rename_table_11 ? io_i_pregs_30 : _GEN_1437; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1439 = 7'h1f == io_i_rename_table_11 ? io_i_pregs_31 : _GEN_1438; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1440 = 7'h20 == io_i_rename_table_11 ? io_i_pregs_32 : _GEN_1439; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1441 = 7'h21 == io_i_rename_table_11 ? io_i_pregs_33 : _GEN_1440; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1442 = 7'h22 == io_i_rename_table_11 ? io_i_pregs_34 : _GEN_1441; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1443 = 7'h23 == io_i_rename_table_11 ? io_i_pregs_35 : _GEN_1442; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1444 = 7'h24 == io_i_rename_table_11 ? io_i_pregs_36 : _GEN_1443; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1445 = 7'h25 == io_i_rename_table_11 ? io_i_pregs_37 : _GEN_1444; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1446 = 7'h26 == io_i_rename_table_11 ? io_i_pregs_38 : _GEN_1445; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1447 = 7'h27 == io_i_rename_table_11 ? io_i_pregs_39 : _GEN_1446; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1448 = 7'h28 == io_i_rename_table_11 ? io_i_pregs_40 : _GEN_1447; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1449 = 7'h29 == io_i_rename_table_11 ? io_i_pregs_41 : _GEN_1448; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1450 = 7'h2a == io_i_rename_table_11 ? io_i_pregs_42 : _GEN_1449; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1451 = 7'h2b == io_i_rename_table_11 ? io_i_pregs_43 : _GEN_1450; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1452 = 7'h2c == io_i_rename_table_11 ? io_i_pregs_44 : _GEN_1451; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1453 = 7'h2d == io_i_rename_table_11 ? io_i_pregs_45 : _GEN_1452; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1454 = 7'h2e == io_i_rename_table_11 ? io_i_pregs_46 : _GEN_1453; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1455 = 7'h2f == io_i_rename_table_11 ? io_i_pregs_47 : _GEN_1454; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1456 = 7'h30 == io_i_rename_table_11 ? io_i_pregs_48 : _GEN_1455; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1457 = 7'h31 == io_i_rename_table_11 ? io_i_pregs_49 : _GEN_1456; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1458 = 7'h32 == io_i_rename_table_11 ? io_i_pregs_50 : _GEN_1457; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1459 = 7'h33 == io_i_rename_table_11 ? io_i_pregs_51 : _GEN_1458; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1460 = 7'h34 == io_i_rename_table_11 ? io_i_pregs_52 : _GEN_1459; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1461 = 7'h35 == io_i_rename_table_11 ? io_i_pregs_53 : _GEN_1460; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1462 = 7'h36 == io_i_rename_table_11 ? io_i_pregs_54 : _GEN_1461; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1463 = 7'h37 == io_i_rename_table_11 ? io_i_pregs_55 : _GEN_1462; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1464 = 7'h38 == io_i_rename_table_11 ? io_i_pregs_56 : _GEN_1463; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1465 = 7'h39 == io_i_rename_table_11 ? io_i_pregs_57 : _GEN_1464; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1466 = 7'h3a == io_i_rename_table_11 ? io_i_pregs_58 : _GEN_1465; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1467 = 7'h3b == io_i_rename_table_11 ? io_i_pregs_59 : _GEN_1466; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1468 = 7'h3c == io_i_rename_table_11 ? io_i_pregs_60 : _GEN_1467; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1469 = 7'h3d == io_i_rename_table_11 ? io_i_pregs_61 : _GEN_1468; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1470 = 7'h3e == io_i_rename_table_11 ? io_i_pregs_62 : _GEN_1469; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1471 = 7'h3f == io_i_rename_table_11 ? io_i_pregs_63 : _GEN_1470; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1472 = 7'h40 == io_i_rename_table_11 ? io_i_pregs_64 : _GEN_1471; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1473 = 7'h41 == io_i_rename_table_11 ? io_i_pregs_65 : _GEN_1472; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1474 = 7'h42 == io_i_rename_table_11 ? io_i_pregs_66 : _GEN_1473; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1475 = 7'h43 == io_i_rename_table_11 ? io_i_pregs_67 : _GEN_1474; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1476 = 7'h44 == io_i_rename_table_11 ? io_i_pregs_68 : _GEN_1475; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1477 = 7'h45 == io_i_rename_table_11 ? io_i_pregs_69 : _GEN_1476; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1478 = 7'h46 == io_i_rename_table_11 ? io_i_pregs_70 : _GEN_1477; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1479 = 7'h47 == io_i_rename_table_11 ? io_i_pregs_71 : _GEN_1478; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1480 = 7'h48 == io_i_rename_table_11 ? io_i_pregs_72 : _GEN_1479; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1481 = 7'h49 == io_i_rename_table_11 ? io_i_pregs_73 : _GEN_1480; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1482 = 7'h4a == io_i_rename_table_11 ? io_i_pregs_74 : _GEN_1481; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1483 = 7'h4b == io_i_rename_table_11 ? io_i_pregs_75 : _GEN_1482; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1484 = 7'h4c == io_i_rename_table_11 ? io_i_pregs_76 : _GEN_1483; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1485 = 7'h4d == io_i_rename_table_11 ? io_i_pregs_77 : _GEN_1484; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1486 = 7'h4e == io_i_rename_table_11 ? io_i_pregs_78 : _GEN_1485; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1487 = 7'h4f == io_i_rename_table_11 ? io_i_pregs_79 : _GEN_1486; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1488 = 7'h50 == io_i_rename_table_11 ? io_i_pregs_80 : _GEN_1487; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1489 = 7'h51 == io_i_rename_table_11 ? io_i_pregs_81 : _GEN_1488; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1490 = 7'h52 == io_i_rename_table_11 ? io_i_pregs_82 : _GEN_1489; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1491 = 7'h53 == io_i_rename_table_11 ? io_i_pregs_83 : _GEN_1490; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1492 = 7'h54 == io_i_rename_table_11 ? io_i_pregs_84 : _GEN_1491; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1493 = 7'h55 == io_i_rename_table_11 ? io_i_pregs_85 : _GEN_1492; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1494 = 7'h56 == io_i_rename_table_11 ? io_i_pregs_86 : _GEN_1493; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1495 = 7'h57 == io_i_rename_table_11 ? io_i_pregs_87 : _GEN_1494; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1496 = 7'h58 == io_i_rename_table_11 ? io_i_pregs_88 : _GEN_1495; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1497 = 7'h59 == io_i_rename_table_11 ? io_i_pregs_89 : _GEN_1496; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1498 = 7'h5a == io_i_rename_table_11 ? io_i_pregs_90 : _GEN_1497; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1499 = 7'h5b == io_i_rename_table_11 ? io_i_pregs_91 : _GEN_1498; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1500 = 7'h5c == io_i_rename_table_11 ? io_i_pregs_92 : _GEN_1499; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1501 = 7'h5d == io_i_rename_table_11 ? io_i_pregs_93 : _GEN_1500; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1502 = 7'h5e == io_i_rename_table_11 ? io_i_pregs_94 : _GEN_1501; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1503 = 7'h5f == io_i_rename_table_11 ? io_i_pregs_95 : _GEN_1502; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1504 = 7'h60 == io_i_rename_table_11 ? io_i_pregs_96 : _GEN_1503; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1505 = 7'h61 == io_i_rename_table_11 ? io_i_pregs_97 : _GEN_1504; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1506 = 7'h62 == io_i_rename_table_11 ? io_i_pregs_98 : _GEN_1505; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1507 = 7'h63 == io_i_rename_table_11 ? io_i_pregs_99 : _GEN_1506; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1508 = 7'h64 == io_i_rename_table_11 ? io_i_pregs_100 : _GEN_1507; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1509 = 7'h65 == io_i_rename_table_11 ? io_i_pregs_101 : _GEN_1508; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1510 = 7'h66 == io_i_rename_table_11 ? io_i_pregs_102 : _GEN_1509; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1511 = 7'h67 == io_i_rename_table_11 ? io_i_pregs_103 : _GEN_1510; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1512 = 7'h68 == io_i_rename_table_11 ? io_i_pregs_104 : _GEN_1511; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1513 = 7'h69 == io_i_rename_table_11 ? io_i_pregs_105 : _GEN_1512; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1514 = 7'h6a == io_i_rename_table_11 ? io_i_pregs_106 : _GEN_1513; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1515 = 7'h6b == io_i_rename_table_11 ? io_i_pregs_107 : _GEN_1514; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1516 = 7'h6c == io_i_rename_table_11 ? io_i_pregs_108 : _GEN_1515; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1517 = 7'h6d == io_i_rename_table_11 ? io_i_pregs_109 : _GEN_1516; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1518 = 7'h6e == io_i_rename_table_11 ? io_i_pregs_110 : _GEN_1517; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1519 = 7'h6f == io_i_rename_table_11 ? io_i_pregs_111 : _GEN_1518; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1520 = 7'h70 == io_i_rename_table_11 ? io_i_pregs_112 : _GEN_1519; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1521 = 7'h71 == io_i_rename_table_11 ? io_i_pregs_113 : _GEN_1520; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1522 = 7'h72 == io_i_rename_table_11 ? io_i_pregs_114 : _GEN_1521; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1523 = 7'h73 == io_i_rename_table_11 ? io_i_pregs_115 : _GEN_1522; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1524 = 7'h74 == io_i_rename_table_11 ? io_i_pregs_116 : _GEN_1523; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1525 = 7'h75 == io_i_rename_table_11 ? io_i_pregs_117 : _GEN_1524; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1526 = 7'h76 == io_i_rename_table_11 ? io_i_pregs_118 : _GEN_1525; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1527 = 7'h77 == io_i_rename_table_11 ? io_i_pregs_119 : _GEN_1526; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1528 = 7'h78 == io_i_rename_table_11 ? io_i_pregs_120 : _GEN_1527; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1529 = 7'h79 == io_i_rename_table_11 ? io_i_pregs_121 : _GEN_1528; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1530 = 7'h7a == io_i_rename_table_11 ? io_i_pregs_122 : _GEN_1529; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1531 = 7'h7b == io_i_rename_table_11 ? io_i_pregs_123 : _GEN_1530; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1532 = 7'h7c == io_i_rename_table_11 ? io_i_pregs_124 : _GEN_1531; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1533 = 7'h7d == io_i_rename_table_11 ? io_i_pregs_125 : _GEN_1532; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1534 = 7'h7e == io_i_rename_table_11 ? io_i_pregs_126 : _GEN_1533; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1537 = 7'h1 == io_i_rename_table_12 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1538 = 7'h2 == io_i_rename_table_12 ? io_i_pregs_2 : _GEN_1537; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1539 = 7'h3 == io_i_rename_table_12 ? io_i_pregs_3 : _GEN_1538; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1540 = 7'h4 == io_i_rename_table_12 ? io_i_pregs_4 : _GEN_1539; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1541 = 7'h5 == io_i_rename_table_12 ? io_i_pregs_5 : _GEN_1540; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1542 = 7'h6 == io_i_rename_table_12 ? io_i_pregs_6 : _GEN_1541; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1543 = 7'h7 == io_i_rename_table_12 ? io_i_pregs_7 : _GEN_1542; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1544 = 7'h8 == io_i_rename_table_12 ? io_i_pregs_8 : _GEN_1543; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1545 = 7'h9 == io_i_rename_table_12 ? io_i_pregs_9 : _GEN_1544; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1546 = 7'ha == io_i_rename_table_12 ? io_i_pregs_10 : _GEN_1545; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1547 = 7'hb == io_i_rename_table_12 ? io_i_pregs_11 : _GEN_1546; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1548 = 7'hc == io_i_rename_table_12 ? io_i_pregs_12 : _GEN_1547; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1549 = 7'hd == io_i_rename_table_12 ? io_i_pregs_13 : _GEN_1548; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1550 = 7'he == io_i_rename_table_12 ? io_i_pregs_14 : _GEN_1549; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1551 = 7'hf == io_i_rename_table_12 ? io_i_pregs_15 : _GEN_1550; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1552 = 7'h10 == io_i_rename_table_12 ? io_i_pregs_16 : _GEN_1551; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1553 = 7'h11 == io_i_rename_table_12 ? io_i_pregs_17 : _GEN_1552; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1554 = 7'h12 == io_i_rename_table_12 ? io_i_pregs_18 : _GEN_1553; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1555 = 7'h13 == io_i_rename_table_12 ? io_i_pregs_19 : _GEN_1554; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1556 = 7'h14 == io_i_rename_table_12 ? io_i_pregs_20 : _GEN_1555; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1557 = 7'h15 == io_i_rename_table_12 ? io_i_pregs_21 : _GEN_1556; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1558 = 7'h16 == io_i_rename_table_12 ? io_i_pregs_22 : _GEN_1557; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1559 = 7'h17 == io_i_rename_table_12 ? io_i_pregs_23 : _GEN_1558; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1560 = 7'h18 == io_i_rename_table_12 ? io_i_pregs_24 : _GEN_1559; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1561 = 7'h19 == io_i_rename_table_12 ? io_i_pregs_25 : _GEN_1560; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1562 = 7'h1a == io_i_rename_table_12 ? io_i_pregs_26 : _GEN_1561; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1563 = 7'h1b == io_i_rename_table_12 ? io_i_pregs_27 : _GEN_1562; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1564 = 7'h1c == io_i_rename_table_12 ? io_i_pregs_28 : _GEN_1563; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1565 = 7'h1d == io_i_rename_table_12 ? io_i_pregs_29 : _GEN_1564; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1566 = 7'h1e == io_i_rename_table_12 ? io_i_pregs_30 : _GEN_1565; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1567 = 7'h1f == io_i_rename_table_12 ? io_i_pregs_31 : _GEN_1566; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1568 = 7'h20 == io_i_rename_table_12 ? io_i_pregs_32 : _GEN_1567; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1569 = 7'h21 == io_i_rename_table_12 ? io_i_pregs_33 : _GEN_1568; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1570 = 7'h22 == io_i_rename_table_12 ? io_i_pregs_34 : _GEN_1569; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1571 = 7'h23 == io_i_rename_table_12 ? io_i_pregs_35 : _GEN_1570; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1572 = 7'h24 == io_i_rename_table_12 ? io_i_pregs_36 : _GEN_1571; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1573 = 7'h25 == io_i_rename_table_12 ? io_i_pregs_37 : _GEN_1572; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1574 = 7'h26 == io_i_rename_table_12 ? io_i_pregs_38 : _GEN_1573; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1575 = 7'h27 == io_i_rename_table_12 ? io_i_pregs_39 : _GEN_1574; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1576 = 7'h28 == io_i_rename_table_12 ? io_i_pregs_40 : _GEN_1575; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1577 = 7'h29 == io_i_rename_table_12 ? io_i_pregs_41 : _GEN_1576; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1578 = 7'h2a == io_i_rename_table_12 ? io_i_pregs_42 : _GEN_1577; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1579 = 7'h2b == io_i_rename_table_12 ? io_i_pregs_43 : _GEN_1578; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1580 = 7'h2c == io_i_rename_table_12 ? io_i_pregs_44 : _GEN_1579; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1581 = 7'h2d == io_i_rename_table_12 ? io_i_pregs_45 : _GEN_1580; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1582 = 7'h2e == io_i_rename_table_12 ? io_i_pregs_46 : _GEN_1581; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1583 = 7'h2f == io_i_rename_table_12 ? io_i_pregs_47 : _GEN_1582; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1584 = 7'h30 == io_i_rename_table_12 ? io_i_pregs_48 : _GEN_1583; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1585 = 7'h31 == io_i_rename_table_12 ? io_i_pregs_49 : _GEN_1584; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1586 = 7'h32 == io_i_rename_table_12 ? io_i_pregs_50 : _GEN_1585; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1587 = 7'h33 == io_i_rename_table_12 ? io_i_pregs_51 : _GEN_1586; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1588 = 7'h34 == io_i_rename_table_12 ? io_i_pregs_52 : _GEN_1587; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1589 = 7'h35 == io_i_rename_table_12 ? io_i_pregs_53 : _GEN_1588; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1590 = 7'h36 == io_i_rename_table_12 ? io_i_pregs_54 : _GEN_1589; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1591 = 7'h37 == io_i_rename_table_12 ? io_i_pregs_55 : _GEN_1590; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1592 = 7'h38 == io_i_rename_table_12 ? io_i_pregs_56 : _GEN_1591; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1593 = 7'h39 == io_i_rename_table_12 ? io_i_pregs_57 : _GEN_1592; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1594 = 7'h3a == io_i_rename_table_12 ? io_i_pregs_58 : _GEN_1593; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1595 = 7'h3b == io_i_rename_table_12 ? io_i_pregs_59 : _GEN_1594; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1596 = 7'h3c == io_i_rename_table_12 ? io_i_pregs_60 : _GEN_1595; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1597 = 7'h3d == io_i_rename_table_12 ? io_i_pregs_61 : _GEN_1596; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1598 = 7'h3e == io_i_rename_table_12 ? io_i_pregs_62 : _GEN_1597; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1599 = 7'h3f == io_i_rename_table_12 ? io_i_pregs_63 : _GEN_1598; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1600 = 7'h40 == io_i_rename_table_12 ? io_i_pregs_64 : _GEN_1599; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1601 = 7'h41 == io_i_rename_table_12 ? io_i_pregs_65 : _GEN_1600; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1602 = 7'h42 == io_i_rename_table_12 ? io_i_pregs_66 : _GEN_1601; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1603 = 7'h43 == io_i_rename_table_12 ? io_i_pregs_67 : _GEN_1602; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1604 = 7'h44 == io_i_rename_table_12 ? io_i_pregs_68 : _GEN_1603; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1605 = 7'h45 == io_i_rename_table_12 ? io_i_pregs_69 : _GEN_1604; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1606 = 7'h46 == io_i_rename_table_12 ? io_i_pregs_70 : _GEN_1605; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1607 = 7'h47 == io_i_rename_table_12 ? io_i_pregs_71 : _GEN_1606; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1608 = 7'h48 == io_i_rename_table_12 ? io_i_pregs_72 : _GEN_1607; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1609 = 7'h49 == io_i_rename_table_12 ? io_i_pregs_73 : _GEN_1608; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1610 = 7'h4a == io_i_rename_table_12 ? io_i_pregs_74 : _GEN_1609; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1611 = 7'h4b == io_i_rename_table_12 ? io_i_pregs_75 : _GEN_1610; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1612 = 7'h4c == io_i_rename_table_12 ? io_i_pregs_76 : _GEN_1611; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1613 = 7'h4d == io_i_rename_table_12 ? io_i_pregs_77 : _GEN_1612; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1614 = 7'h4e == io_i_rename_table_12 ? io_i_pregs_78 : _GEN_1613; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1615 = 7'h4f == io_i_rename_table_12 ? io_i_pregs_79 : _GEN_1614; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1616 = 7'h50 == io_i_rename_table_12 ? io_i_pregs_80 : _GEN_1615; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1617 = 7'h51 == io_i_rename_table_12 ? io_i_pregs_81 : _GEN_1616; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1618 = 7'h52 == io_i_rename_table_12 ? io_i_pregs_82 : _GEN_1617; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1619 = 7'h53 == io_i_rename_table_12 ? io_i_pregs_83 : _GEN_1618; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1620 = 7'h54 == io_i_rename_table_12 ? io_i_pregs_84 : _GEN_1619; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1621 = 7'h55 == io_i_rename_table_12 ? io_i_pregs_85 : _GEN_1620; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1622 = 7'h56 == io_i_rename_table_12 ? io_i_pregs_86 : _GEN_1621; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1623 = 7'h57 == io_i_rename_table_12 ? io_i_pregs_87 : _GEN_1622; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1624 = 7'h58 == io_i_rename_table_12 ? io_i_pregs_88 : _GEN_1623; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1625 = 7'h59 == io_i_rename_table_12 ? io_i_pregs_89 : _GEN_1624; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1626 = 7'h5a == io_i_rename_table_12 ? io_i_pregs_90 : _GEN_1625; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1627 = 7'h5b == io_i_rename_table_12 ? io_i_pregs_91 : _GEN_1626; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1628 = 7'h5c == io_i_rename_table_12 ? io_i_pregs_92 : _GEN_1627; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1629 = 7'h5d == io_i_rename_table_12 ? io_i_pregs_93 : _GEN_1628; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1630 = 7'h5e == io_i_rename_table_12 ? io_i_pregs_94 : _GEN_1629; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1631 = 7'h5f == io_i_rename_table_12 ? io_i_pregs_95 : _GEN_1630; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1632 = 7'h60 == io_i_rename_table_12 ? io_i_pregs_96 : _GEN_1631; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1633 = 7'h61 == io_i_rename_table_12 ? io_i_pregs_97 : _GEN_1632; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1634 = 7'h62 == io_i_rename_table_12 ? io_i_pregs_98 : _GEN_1633; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1635 = 7'h63 == io_i_rename_table_12 ? io_i_pregs_99 : _GEN_1634; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1636 = 7'h64 == io_i_rename_table_12 ? io_i_pregs_100 : _GEN_1635; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1637 = 7'h65 == io_i_rename_table_12 ? io_i_pregs_101 : _GEN_1636; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1638 = 7'h66 == io_i_rename_table_12 ? io_i_pregs_102 : _GEN_1637; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1639 = 7'h67 == io_i_rename_table_12 ? io_i_pregs_103 : _GEN_1638; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1640 = 7'h68 == io_i_rename_table_12 ? io_i_pregs_104 : _GEN_1639; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1641 = 7'h69 == io_i_rename_table_12 ? io_i_pregs_105 : _GEN_1640; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1642 = 7'h6a == io_i_rename_table_12 ? io_i_pregs_106 : _GEN_1641; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1643 = 7'h6b == io_i_rename_table_12 ? io_i_pregs_107 : _GEN_1642; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1644 = 7'h6c == io_i_rename_table_12 ? io_i_pregs_108 : _GEN_1643; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1645 = 7'h6d == io_i_rename_table_12 ? io_i_pregs_109 : _GEN_1644; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1646 = 7'h6e == io_i_rename_table_12 ? io_i_pregs_110 : _GEN_1645; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1647 = 7'h6f == io_i_rename_table_12 ? io_i_pregs_111 : _GEN_1646; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1648 = 7'h70 == io_i_rename_table_12 ? io_i_pregs_112 : _GEN_1647; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1649 = 7'h71 == io_i_rename_table_12 ? io_i_pregs_113 : _GEN_1648; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1650 = 7'h72 == io_i_rename_table_12 ? io_i_pregs_114 : _GEN_1649; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1651 = 7'h73 == io_i_rename_table_12 ? io_i_pregs_115 : _GEN_1650; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1652 = 7'h74 == io_i_rename_table_12 ? io_i_pregs_116 : _GEN_1651; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1653 = 7'h75 == io_i_rename_table_12 ? io_i_pregs_117 : _GEN_1652; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1654 = 7'h76 == io_i_rename_table_12 ? io_i_pregs_118 : _GEN_1653; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1655 = 7'h77 == io_i_rename_table_12 ? io_i_pregs_119 : _GEN_1654; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1656 = 7'h78 == io_i_rename_table_12 ? io_i_pregs_120 : _GEN_1655; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1657 = 7'h79 == io_i_rename_table_12 ? io_i_pregs_121 : _GEN_1656; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1658 = 7'h7a == io_i_rename_table_12 ? io_i_pregs_122 : _GEN_1657; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1659 = 7'h7b == io_i_rename_table_12 ? io_i_pregs_123 : _GEN_1658; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1660 = 7'h7c == io_i_rename_table_12 ? io_i_pregs_124 : _GEN_1659; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1661 = 7'h7d == io_i_rename_table_12 ? io_i_pregs_125 : _GEN_1660; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1662 = 7'h7e == io_i_rename_table_12 ? io_i_pregs_126 : _GEN_1661; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1665 = 7'h1 == io_i_rename_table_13 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1666 = 7'h2 == io_i_rename_table_13 ? io_i_pregs_2 : _GEN_1665; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1667 = 7'h3 == io_i_rename_table_13 ? io_i_pregs_3 : _GEN_1666; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1668 = 7'h4 == io_i_rename_table_13 ? io_i_pregs_4 : _GEN_1667; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1669 = 7'h5 == io_i_rename_table_13 ? io_i_pregs_5 : _GEN_1668; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1670 = 7'h6 == io_i_rename_table_13 ? io_i_pregs_6 : _GEN_1669; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1671 = 7'h7 == io_i_rename_table_13 ? io_i_pregs_7 : _GEN_1670; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1672 = 7'h8 == io_i_rename_table_13 ? io_i_pregs_8 : _GEN_1671; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1673 = 7'h9 == io_i_rename_table_13 ? io_i_pregs_9 : _GEN_1672; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1674 = 7'ha == io_i_rename_table_13 ? io_i_pregs_10 : _GEN_1673; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1675 = 7'hb == io_i_rename_table_13 ? io_i_pregs_11 : _GEN_1674; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1676 = 7'hc == io_i_rename_table_13 ? io_i_pregs_12 : _GEN_1675; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1677 = 7'hd == io_i_rename_table_13 ? io_i_pregs_13 : _GEN_1676; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1678 = 7'he == io_i_rename_table_13 ? io_i_pregs_14 : _GEN_1677; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1679 = 7'hf == io_i_rename_table_13 ? io_i_pregs_15 : _GEN_1678; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1680 = 7'h10 == io_i_rename_table_13 ? io_i_pregs_16 : _GEN_1679; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1681 = 7'h11 == io_i_rename_table_13 ? io_i_pregs_17 : _GEN_1680; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1682 = 7'h12 == io_i_rename_table_13 ? io_i_pregs_18 : _GEN_1681; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1683 = 7'h13 == io_i_rename_table_13 ? io_i_pregs_19 : _GEN_1682; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1684 = 7'h14 == io_i_rename_table_13 ? io_i_pregs_20 : _GEN_1683; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1685 = 7'h15 == io_i_rename_table_13 ? io_i_pregs_21 : _GEN_1684; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1686 = 7'h16 == io_i_rename_table_13 ? io_i_pregs_22 : _GEN_1685; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1687 = 7'h17 == io_i_rename_table_13 ? io_i_pregs_23 : _GEN_1686; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1688 = 7'h18 == io_i_rename_table_13 ? io_i_pregs_24 : _GEN_1687; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1689 = 7'h19 == io_i_rename_table_13 ? io_i_pregs_25 : _GEN_1688; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1690 = 7'h1a == io_i_rename_table_13 ? io_i_pregs_26 : _GEN_1689; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1691 = 7'h1b == io_i_rename_table_13 ? io_i_pregs_27 : _GEN_1690; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1692 = 7'h1c == io_i_rename_table_13 ? io_i_pregs_28 : _GEN_1691; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1693 = 7'h1d == io_i_rename_table_13 ? io_i_pregs_29 : _GEN_1692; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1694 = 7'h1e == io_i_rename_table_13 ? io_i_pregs_30 : _GEN_1693; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1695 = 7'h1f == io_i_rename_table_13 ? io_i_pregs_31 : _GEN_1694; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1696 = 7'h20 == io_i_rename_table_13 ? io_i_pregs_32 : _GEN_1695; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1697 = 7'h21 == io_i_rename_table_13 ? io_i_pregs_33 : _GEN_1696; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1698 = 7'h22 == io_i_rename_table_13 ? io_i_pregs_34 : _GEN_1697; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1699 = 7'h23 == io_i_rename_table_13 ? io_i_pregs_35 : _GEN_1698; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1700 = 7'h24 == io_i_rename_table_13 ? io_i_pregs_36 : _GEN_1699; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1701 = 7'h25 == io_i_rename_table_13 ? io_i_pregs_37 : _GEN_1700; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1702 = 7'h26 == io_i_rename_table_13 ? io_i_pregs_38 : _GEN_1701; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1703 = 7'h27 == io_i_rename_table_13 ? io_i_pregs_39 : _GEN_1702; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1704 = 7'h28 == io_i_rename_table_13 ? io_i_pregs_40 : _GEN_1703; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1705 = 7'h29 == io_i_rename_table_13 ? io_i_pregs_41 : _GEN_1704; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1706 = 7'h2a == io_i_rename_table_13 ? io_i_pregs_42 : _GEN_1705; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1707 = 7'h2b == io_i_rename_table_13 ? io_i_pregs_43 : _GEN_1706; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1708 = 7'h2c == io_i_rename_table_13 ? io_i_pregs_44 : _GEN_1707; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1709 = 7'h2d == io_i_rename_table_13 ? io_i_pregs_45 : _GEN_1708; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1710 = 7'h2e == io_i_rename_table_13 ? io_i_pregs_46 : _GEN_1709; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1711 = 7'h2f == io_i_rename_table_13 ? io_i_pregs_47 : _GEN_1710; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1712 = 7'h30 == io_i_rename_table_13 ? io_i_pregs_48 : _GEN_1711; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1713 = 7'h31 == io_i_rename_table_13 ? io_i_pregs_49 : _GEN_1712; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1714 = 7'h32 == io_i_rename_table_13 ? io_i_pregs_50 : _GEN_1713; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1715 = 7'h33 == io_i_rename_table_13 ? io_i_pregs_51 : _GEN_1714; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1716 = 7'h34 == io_i_rename_table_13 ? io_i_pregs_52 : _GEN_1715; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1717 = 7'h35 == io_i_rename_table_13 ? io_i_pregs_53 : _GEN_1716; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1718 = 7'h36 == io_i_rename_table_13 ? io_i_pregs_54 : _GEN_1717; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1719 = 7'h37 == io_i_rename_table_13 ? io_i_pregs_55 : _GEN_1718; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1720 = 7'h38 == io_i_rename_table_13 ? io_i_pregs_56 : _GEN_1719; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1721 = 7'h39 == io_i_rename_table_13 ? io_i_pregs_57 : _GEN_1720; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1722 = 7'h3a == io_i_rename_table_13 ? io_i_pregs_58 : _GEN_1721; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1723 = 7'h3b == io_i_rename_table_13 ? io_i_pregs_59 : _GEN_1722; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1724 = 7'h3c == io_i_rename_table_13 ? io_i_pregs_60 : _GEN_1723; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1725 = 7'h3d == io_i_rename_table_13 ? io_i_pregs_61 : _GEN_1724; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1726 = 7'h3e == io_i_rename_table_13 ? io_i_pregs_62 : _GEN_1725; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1727 = 7'h3f == io_i_rename_table_13 ? io_i_pregs_63 : _GEN_1726; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1728 = 7'h40 == io_i_rename_table_13 ? io_i_pregs_64 : _GEN_1727; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1729 = 7'h41 == io_i_rename_table_13 ? io_i_pregs_65 : _GEN_1728; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1730 = 7'h42 == io_i_rename_table_13 ? io_i_pregs_66 : _GEN_1729; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1731 = 7'h43 == io_i_rename_table_13 ? io_i_pregs_67 : _GEN_1730; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1732 = 7'h44 == io_i_rename_table_13 ? io_i_pregs_68 : _GEN_1731; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1733 = 7'h45 == io_i_rename_table_13 ? io_i_pregs_69 : _GEN_1732; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1734 = 7'h46 == io_i_rename_table_13 ? io_i_pregs_70 : _GEN_1733; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1735 = 7'h47 == io_i_rename_table_13 ? io_i_pregs_71 : _GEN_1734; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1736 = 7'h48 == io_i_rename_table_13 ? io_i_pregs_72 : _GEN_1735; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1737 = 7'h49 == io_i_rename_table_13 ? io_i_pregs_73 : _GEN_1736; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1738 = 7'h4a == io_i_rename_table_13 ? io_i_pregs_74 : _GEN_1737; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1739 = 7'h4b == io_i_rename_table_13 ? io_i_pregs_75 : _GEN_1738; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1740 = 7'h4c == io_i_rename_table_13 ? io_i_pregs_76 : _GEN_1739; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1741 = 7'h4d == io_i_rename_table_13 ? io_i_pregs_77 : _GEN_1740; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1742 = 7'h4e == io_i_rename_table_13 ? io_i_pregs_78 : _GEN_1741; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1743 = 7'h4f == io_i_rename_table_13 ? io_i_pregs_79 : _GEN_1742; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1744 = 7'h50 == io_i_rename_table_13 ? io_i_pregs_80 : _GEN_1743; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1745 = 7'h51 == io_i_rename_table_13 ? io_i_pregs_81 : _GEN_1744; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1746 = 7'h52 == io_i_rename_table_13 ? io_i_pregs_82 : _GEN_1745; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1747 = 7'h53 == io_i_rename_table_13 ? io_i_pregs_83 : _GEN_1746; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1748 = 7'h54 == io_i_rename_table_13 ? io_i_pregs_84 : _GEN_1747; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1749 = 7'h55 == io_i_rename_table_13 ? io_i_pregs_85 : _GEN_1748; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1750 = 7'h56 == io_i_rename_table_13 ? io_i_pregs_86 : _GEN_1749; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1751 = 7'h57 == io_i_rename_table_13 ? io_i_pregs_87 : _GEN_1750; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1752 = 7'h58 == io_i_rename_table_13 ? io_i_pregs_88 : _GEN_1751; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1753 = 7'h59 == io_i_rename_table_13 ? io_i_pregs_89 : _GEN_1752; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1754 = 7'h5a == io_i_rename_table_13 ? io_i_pregs_90 : _GEN_1753; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1755 = 7'h5b == io_i_rename_table_13 ? io_i_pregs_91 : _GEN_1754; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1756 = 7'h5c == io_i_rename_table_13 ? io_i_pregs_92 : _GEN_1755; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1757 = 7'h5d == io_i_rename_table_13 ? io_i_pregs_93 : _GEN_1756; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1758 = 7'h5e == io_i_rename_table_13 ? io_i_pregs_94 : _GEN_1757; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1759 = 7'h5f == io_i_rename_table_13 ? io_i_pregs_95 : _GEN_1758; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1760 = 7'h60 == io_i_rename_table_13 ? io_i_pregs_96 : _GEN_1759; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1761 = 7'h61 == io_i_rename_table_13 ? io_i_pregs_97 : _GEN_1760; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1762 = 7'h62 == io_i_rename_table_13 ? io_i_pregs_98 : _GEN_1761; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1763 = 7'h63 == io_i_rename_table_13 ? io_i_pregs_99 : _GEN_1762; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1764 = 7'h64 == io_i_rename_table_13 ? io_i_pregs_100 : _GEN_1763; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1765 = 7'h65 == io_i_rename_table_13 ? io_i_pregs_101 : _GEN_1764; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1766 = 7'h66 == io_i_rename_table_13 ? io_i_pregs_102 : _GEN_1765; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1767 = 7'h67 == io_i_rename_table_13 ? io_i_pregs_103 : _GEN_1766; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1768 = 7'h68 == io_i_rename_table_13 ? io_i_pregs_104 : _GEN_1767; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1769 = 7'h69 == io_i_rename_table_13 ? io_i_pregs_105 : _GEN_1768; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1770 = 7'h6a == io_i_rename_table_13 ? io_i_pregs_106 : _GEN_1769; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1771 = 7'h6b == io_i_rename_table_13 ? io_i_pregs_107 : _GEN_1770; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1772 = 7'h6c == io_i_rename_table_13 ? io_i_pregs_108 : _GEN_1771; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1773 = 7'h6d == io_i_rename_table_13 ? io_i_pregs_109 : _GEN_1772; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1774 = 7'h6e == io_i_rename_table_13 ? io_i_pregs_110 : _GEN_1773; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1775 = 7'h6f == io_i_rename_table_13 ? io_i_pregs_111 : _GEN_1774; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1776 = 7'h70 == io_i_rename_table_13 ? io_i_pregs_112 : _GEN_1775; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1777 = 7'h71 == io_i_rename_table_13 ? io_i_pregs_113 : _GEN_1776; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1778 = 7'h72 == io_i_rename_table_13 ? io_i_pregs_114 : _GEN_1777; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1779 = 7'h73 == io_i_rename_table_13 ? io_i_pregs_115 : _GEN_1778; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1780 = 7'h74 == io_i_rename_table_13 ? io_i_pregs_116 : _GEN_1779; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1781 = 7'h75 == io_i_rename_table_13 ? io_i_pregs_117 : _GEN_1780; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1782 = 7'h76 == io_i_rename_table_13 ? io_i_pregs_118 : _GEN_1781; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1783 = 7'h77 == io_i_rename_table_13 ? io_i_pregs_119 : _GEN_1782; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1784 = 7'h78 == io_i_rename_table_13 ? io_i_pregs_120 : _GEN_1783; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1785 = 7'h79 == io_i_rename_table_13 ? io_i_pregs_121 : _GEN_1784; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1786 = 7'h7a == io_i_rename_table_13 ? io_i_pregs_122 : _GEN_1785; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1787 = 7'h7b == io_i_rename_table_13 ? io_i_pregs_123 : _GEN_1786; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1788 = 7'h7c == io_i_rename_table_13 ? io_i_pregs_124 : _GEN_1787; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1789 = 7'h7d == io_i_rename_table_13 ? io_i_pregs_125 : _GEN_1788; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1790 = 7'h7e == io_i_rename_table_13 ? io_i_pregs_126 : _GEN_1789; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1793 = 7'h1 == io_i_rename_table_14 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1794 = 7'h2 == io_i_rename_table_14 ? io_i_pregs_2 : _GEN_1793; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1795 = 7'h3 == io_i_rename_table_14 ? io_i_pregs_3 : _GEN_1794; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1796 = 7'h4 == io_i_rename_table_14 ? io_i_pregs_4 : _GEN_1795; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1797 = 7'h5 == io_i_rename_table_14 ? io_i_pregs_5 : _GEN_1796; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1798 = 7'h6 == io_i_rename_table_14 ? io_i_pregs_6 : _GEN_1797; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1799 = 7'h7 == io_i_rename_table_14 ? io_i_pregs_7 : _GEN_1798; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1800 = 7'h8 == io_i_rename_table_14 ? io_i_pregs_8 : _GEN_1799; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1801 = 7'h9 == io_i_rename_table_14 ? io_i_pregs_9 : _GEN_1800; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1802 = 7'ha == io_i_rename_table_14 ? io_i_pregs_10 : _GEN_1801; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1803 = 7'hb == io_i_rename_table_14 ? io_i_pregs_11 : _GEN_1802; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1804 = 7'hc == io_i_rename_table_14 ? io_i_pregs_12 : _GEN_1803; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1805 = 7'hd == io_i_rename_table_14 ? io_i_pregs_13 : _GEN_1804; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1806 = 7'he == io_i_rename_table_14 ? io_i_pregs_14 : _GEN_1805; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1807 = 7'hf == io_i_rename_table_14 ? io_i_pregs_15 : _GEN_1806; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1808 = 7'h10 == io_i_rename_table_14 ? io_i_pregs_16 : _GEN_1807; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1809 = 7'h11 == io_i_rename_table_14 ? io_i_pregs_17 : _GEN_1808; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1810 = 7'h12 == io_i_rename_table_14 ? io_i_pregs_18 : _GEN_1809; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1811 = 7'h13 == io_i_rename_table_14 ? io_i_pregs_19 : _GEN_1810; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1812 = 7'h14 == io_i_rename_table_14 ? io_i_pregs_20 : _GEN_1811; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1813 = 7'h15 == io_i_rename_table_14 ? io_i_pregs_21 : _GEN_1812; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1814 = 7'h16 == io_i_rename_table_14 ? io_i_pregs_22 : _GEN_1813; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1815 = 7'h17 == io_i_rename_table_14 ? io_i_pregs_23 : _GEN_1814; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1816 = 7'h18 == io_i_rename_table_14 ? io_i_pregs_24 : _GEN_1815; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1817 = 7'h19 == io_i_rename_table_14 ? io_i_pregs_25 : _GEN_1816; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1818 = 7'h1a == io_i_rename_table_14 ? io_i_pregs_26 : _GEN_1817; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1819 = 7'h1b == io_i_rename_table_14 ? io_i_pregs_27 : _GEN_1818; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1820 = 7'h1c == io_i_rename_table_14 ? io_i_pregs_28 : _GEN_1819; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1821 = 7'h1d == io_i_rename_table_14 ? io_i_pregs_29 : _GEN_1820; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1822 = 7'h1e == io_i_rename_table_14 ? io_i_pregs_30 : _GEN_1821; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1823 = 7'h1f == io_i_rename_table_14 ? io_i_pregs_31 : _GEN_1822; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1824 = 7'h20 == io_i_rename_table_14 ? io_i_pregs_32 : _GEN_1823; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1825 = 7'h21 == io_i_rename_table_14 ? io_i_pregs_33 : _GEN_1824; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1826 = 7'h22 == io_i_rename_table_14 ? io_i_pregs_34 : _GEN_1825; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1827 = 7'h23 == io_i_rename_table_14 ? io_i_pregs_35 : _GEN_1826; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1828 = 7'h24 == io_i_rename_table_14 ? io_i_pregs_36 : _GEN_1827; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1829 = 7'h25 == io_i_rename_table_14 ? io_i_pregs_37 : _GEN_1828; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1830 = 7'h26 == io_i_rename_table_14 ? io_i_pregs_38 : _GEN_1829; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1831 = 7'h27 == io_i_rename_table_14 ? io_i_pregs_39 : _GEN_1830; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1832 = 7'h28 == io_i_rename_table_14 ? io_i_pregs_40 : _GEN_1831; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1833 = 7'h29 == io_i_rename_table_14 ? io_i_pregs_41 : _GEN_1832; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1834 = 7'h2a == io_i_rename_table_14 ? io_i_pregs_42 : _GEN_1833; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1835 = 7'h2b == io_i_rename_table_14 ? io_i_pregs_43 : _GEN_1834; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1836 = 7'h2c == io_i_rename_table_14 ? io_i_pregs_44 : _GEN_1835; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1837 = 7'h2d == io_i_rename_table_14 ? io_i_pregs_45 : _GEN_1836; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1838 = 7'h2e == io_i_rename_table_14 ? io_i_pregs_46 : _GEN_1837; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1839 = 7'h2f == io_i_rename_table_14 ? io_i_pregs_47 : _GEN_1838; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1840 = 7'h30 == io_i_rename_table_14 ? io_i_pregs_48 : _GEN_1839; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1841 = 7'h31 == io_i_rename_table_14 ? io_i_pregs_49 : _GEN_1840; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1842 = 7'h32 == io_i_rename_table_14 ? io_i_pregs_50 : _GEN_1841; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1843 = 7'h33 == io_i_rename_table_14 ? io_i_pregs_51 : _GEN_1842; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1844 = 7'h34 == io_i_rename_table_14 ? io_i_pregs_52 : _GEN_1843; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1845 = 7'h35 == io_i_rename_table_14 ? io_i_pregs_53 : _GEN_1844; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1846 = 7'h36 == io_i_rename_table_14 ? io_i_pregs_54 : _GEN_1845; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1847 = 7'h37 == io_i_rename_table_14 ? io_i_pregs_55 : _GEN_1846; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1848 = 7'h38 == io_i_rename_table_14 ? io_i_pregs_56 : _GEN_1847; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1849 = 7'h39 == io_i_rename_table_14 ? io_i_pregs_57 : _GEN_1848; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1850 = 7'h3a == io_i_rename_table_14 ? io_i_pregs_58 : _GEN_1849; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1851 = 7'h3b == io_i_rename_table_14 ? io_i_pregs_59 : _GEN_1850; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1852 = 7'h3c == io_i_rename_table_14 ? io_i_pregs_60 : _GEN_1851; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1853 = 7'h3d == io_i_rename_table_14 ? io_i_pregs_61 : _GEN_1852; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1854 = 7'h3e == io_i_rename_table_14 ? io_i_pregs_62 : _GEN_1853; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1855 = 7'h3f == io_i_rename_table_14 ? io_i_pregs_63 : _GEN_1854; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1856 = 7'h40 == io_i_rename_table_14 ? io_i_pregs_64 : _GEN_1855; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1857 = 7'h41 == io_i_rename_table_14 ? io_i_pregs_65 : _GEN_1856; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1858 = 7'h42 == io_i_rename_table_14 ? io_i_pregs_66 : _GEN_1857; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1859 = 7'h43 == io_i_rename_table_14 ? io_i_pregs_67 : _GEN_1858; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1860 = 7'h44 == io_i_rename_table_14 ? io_i_pregs_68 : _GEN_1859; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1861 = 7'h45 == io_i_rename_table_14 ? io_i_pregs_69 : _GEN_1860; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1862 = 7'h46 == io_i_rename_table_14 ? io_i_pregs_70 : _GEN_1861; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1863 = 7'h47 == io_i_rename_table_14 ? io_i_pregs_71 : _GEN_1862; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1864 = 7'h48 == io_i_rename_table_14 ? io_i_pregs_72 : _GEN_1863; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1865 = 7'h49 == io_i_rename_table_14 ? io_i_pregs_73 : _GEN_1864; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1866 = 7'h4a == io_i_rename_table_14 ? io_i_pregs_74 : _GEN_1865; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1867 = 7'h4b == io_i_rename_table_14 ? io_i_pregs_75 : _GEN_1866; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1868 = 7'h4c == io_i_rename_table_14 ? io_i_pregs_76 : _GEN_1867; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1869 = 7'h4d == io_i_rename_table_14 ? io_i_pregs_77 : _GEN_1868; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1870 = 7'h4e == io_i_rename_table_14 ? io_i_pregs_78 : _GEN_1869; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1871 = 7'h4f == io_i_rename_table_14 ? io_i_pregs_79 : _GEN_1870; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1872 = 7'h50 == io_i_rename_table_14 ? io_i_pregs_80 : _GEN_1871; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1873 = 7'h51 == io_i_rename_table_14 ? io_i_pregs_81 : _GEN_1872; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1874 = 7'h52 == io_i_rename_table_14 ? io_i_pregs_82 : _GEN_1873; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1875 = 7'h53 == io_i_rename_table_14 ? io_i_pregs_83 : _GEN_1874; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1876 = 7'h54 == io_i_rename_table_14 ? io_i_pregs_84 : _GEN_1875; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1877 = 7'h55 == io_i_rename_table_14 ? io_i_pregs_85 : _GEN_1876; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1878 = 7'h56 == io_i_rename_table_14 ? io_i_pregs_86 : _GEN_1877; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1879 = 7'h57 == io_i_rename_table_14 ? io_i_pregs_87 : _GEN_1878; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1880 = 7'h58 == io_i_rename_table_14 ? io_i_pregs_88 : _GEN_1879; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1881 = 7'h59 == io_i_rename_table_14 ? io_i_pregs_89 : _GEN_1880; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1882 = 7'h5a == io_i_rename_table_14 ? io_i_pregs_90 : _GEN_1881; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1883 = 7'h5b == io_i_rename_table_14 ? io_i_pregs_91 : _GEN_1882; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1884 = 7'h5c == io_i_rename_table_14 ? io_i_pregs_92 : _GEN_1883; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1885 = 7'h5d == io_i_rename_table_14 ? io_i_pregs_93 : _GEN_1884; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1886 = 7'h5e == io_i_rename_table_14 ? io_i_pregs_94 : _GEN_1885; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1887 = 7'h5f == io_i_rename_table_14 ? io_i_pregs_95 : _GEN_1886; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1888 = 7'h60 == io_i_rename_table_14 ? io_i_pregs_96 : _GEN_1887; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1889 = 7'h61 == io_i_rename_table_14 ? io_i_pregs_97 : _GEN_1888; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1890 = 7'h62 == io_i_rename_table_14 ? io_i_pregs_98 : _GEN_1889; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1891 = 7'h63 == io_i_rename_table_14 ? io_i_pregs_99 : _GEN_1890; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1892 = 7'h64 == io_i_rename_table_14 ? io_i_pregs_100 : _GEN_1891; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1893 = 7'h65 == io_i_rename_table_14 ? io_i_pregs_101 : _GEN_1892; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1894 = 7'h66 == io_i_rename_table_14 ? io_i_pregs_102 : _GEN_1893; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1895 = 7'h67 == io_i_rename_table_14 ? io_i_pregs_103 : _GEN_1894; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1896 = 7'h68 == io_i_rename_table_14 ? io_i_pregs_104 : _GEN_1895; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1897 = 7'h69 == io_i_rename_table_14 ? io_i_pregs_105 : _GEN_1896; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1898 = 7'h6a == io_i_rename_table_14 ? io_i_pregs_106 : _GEN_1897; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1899 = 7'h6b == io_i_rename_table_14 ? io_i_pregs_107 : _GEN_1898; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1900 = 7'h6c == io_i_rename_table_14 ? io_i_pregs_108 : _GEN_1899; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1901 = 7'h6d == io_i_rename_table_14 ? io_i_pregs_109 : _GEN_1900; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1902 = 7'h6e == io_i_rename_table_14 ? io_i_pregs_110 : _GEN_1901; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1903 = 7'h6f == io_i_rename_table_14 ? io_i_pregs_111 : _GEN_1902; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1904 = 7'h70 == io_i_rename_table_14 ? io_i_pregs_112 : _GEN_1903; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1905 = 7'h71 == io_i_rename_table_14 ? io_i_pregs_113 : _GEN_1904; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1906 = 7'h72 == io_i_rename_table_14 ? io_i_pregs_114 : _GEN_1905; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1907 = 7'h73 == io_i_rename_table_14 ? io_i_pregs_115 : _GEN_1906; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1908 = 7'h74 == io_i_rename_table_14 ? io_i_pregs_116 : _GEN_1907; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1909 = 7'h75 == io_i_rename_table_14 ? io_i_pregs_117 : _GEN_1908; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1910 = 7'h76 == io_i_rename_table_14 ? io_i_pregs_118 : _GEN_1909; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1911 = 7'h77 == io_i_rename_table_14 ? io_i_pregs_119 : _GEN_1910; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1912 = 7'h78 == io_i_rename_table_14 ? io_i_pregs_120 : _GEN_1911; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1913 = 7'h79 == io_i_rename_table_14 ? io_i_pregs_121 : _GEN_1912; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1914 = 7'h7a == io_i_rename_table_14 ? io_i_pregs_122 : _GEN_1913; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1915 = 7'h7b == io_i_rename_table_14 ? io_i_pregs_123 : _GEN_1914; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1916 = 7'h7c == io_i_rename_table_14 ? io_i_pregs_124 : _GEN_1915; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1917 = 7'h7d == io_i_rename_table_14 ? io_i_pregs_125 : _GEN_1916; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1918 = 7'h7e == io_i_rename_table_14 ? io_i_pregs_126 : _GEN_1917; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1921 = 7'h1 == io_i_rename_table_15 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1922 = 7'h2 == io_i_rename_table_15 ? io_i_pregs_2 : _GEN_1921; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1923 = 7'h3 == io_i_rename_table_15 ? io_i_pregs_3 : _GEN_1922; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1924 = 7'h4 == io_i_rename_table_15 ? io_i_pregs_4 : _GEN_1923; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1925 = 7'h5 == io_i_rename_table_15 ? io_i_pregs_5 : _GEN_1924; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1926 = 7'h6 == io_i_rename_table_15 ? io_i_pregs_6 : _GEN_1925; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1927 = 7'h7 == io_i_rename_table_15 ? io_i_pregs_7 : _GEN_1926; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1928 = 7'h8 == io_i_rename_table_15 ? io_i_pregs_8 : _GEN_1927; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1929 = 7'h9 == io_i_rename_table_15 ? io_i_pregs_9 : _GEN_1928; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1930 = 7'ha == io_i_rename_table_15 ? io_i_pregs_10 : _GEN_1929; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1931 = 7'hb == io_i_rename_table_15 ? io_i_pregs_11 : _GEN_1930; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1932 = 7'hc == io_i_rename_table_15 ? io_i_pregs_12 : _GEN_1931; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1933 = 7'hd == io_i_rename_table_15 ? io_i_pregs_13 : _GEN_1932; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1934 = 7'he == io_i_rename_table_15 ? io_i_pregs_14 : _GEN_1933; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1935 = 7'hf == io_i_rename_table_15 ? io_i_pregs_15 : _GEN_1934; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1936 = 7'h10 == io_i_rename_table_15 ? io_i_pregs_16 : _GEN_1935; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1937 = 7'h11 == io_i_rename_table_15 ? io_i_pregs_17 : _GEN_1936; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1938 = 7'h12 == io_i_rename_table_15 ? io_i_pregs_18 : _GEN_1937; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1939 = 7'h13 == io_i_rename_table_15 ? io_i_pregs_19 : _GEN_1938; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1940 = 7'h14 == io_i_rename_table_15 ? io_i_pregs_20 : _GEN_1939; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1941 = 7'h15 == io_i_rename_table_15 ? io_i_pregs_21 : _GEN_1940; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1942 = 7'h16 == io_i_rename_table_15 ? io_i_pregs_22 : _GEN_1941; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1943 = 7'h17 == io_i_rename_table_15 ? io_i_pregs_23 : _GEN_1942; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1944 = 7'h18 == io_i_rename_table_15 ? io_i_pregs_24 : _GEN_1943; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1945 = 7'h19 == io_i_rename_table_15 ? io_i_pregs_25 : _GEN_1944; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1946 = 7'h1a == io_i_rename_table_15 ? io_i_pregs_26 : _GEN_1945; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1947 = 7'h1b == io_i_rename_table_15 ? io_i_pregs_27 : _GEN_1946; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1948 = 7'h1c == io_i_rename_table_15 ? io_i_pregs_28 : _GEN_1947; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1949 = 7'h1d == io_i_rename_table_15 ? io_i_pregs_29 : _GEN_1948; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1950 = 7'h1e == io_i_rename_table_15 ? io_i_pregs_30 : _GEN_1949; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1951 = 7'h1f == io_i_rename_table_15 ? io_i_pregs_31 : _GEN_1950; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1952 = 7'h20 == io_i_rename_table_15 ? io_i_pregs_32 : _GEN_1951; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1953 = 7'h21 == io_i_rename_table_15 ? io_i_pregs_33 : _GEN_1952; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1954 = 7'h22 == io_i_rename_table_15 ? io_i_pregs_34 : _GEN_1953; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1955 = 7'h23 == io_i_rename_table_15 ? io_i_pregs_35 : _GEN_1954; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1956 = 7'h24 == io_i_rename_table_15 ? io_i_pregs_36 : _GEN_1955; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1957 = 7'h25 == io_i_rename_table_15 ? io_i_pregs_37 : _GEN_1956; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1958 = 7'h26 == io_i_rename_table_15 ? io_i_pregs_38 : _GEN_1957; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1959 = 7'h27 == io_i_rename_table_15 ? io_i_pregs_39 : _GEN_1958; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1960 = 7'h28 == io_i_rename_table_15 ? io_i_pregs_40 : _GEN_1959; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1961 = 7'h29 == io_i_rename_table_15 ? io_i_pregs_41 : _GEN_1960; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1962 = 7'h2a == io_i_rename_table_15 ? io_i_pregs_42 : _GEN_1961; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1963 = 7'h2b == io_i_rename_table_15 ? io_i_pregs_43 : _GEN_1962; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1964 = 7'h2c == io_i_rename_table_15 ? io_i_pregs_44 : _GEN_1963; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1965 = 7'h2d == io_i_rename_table_15 ? io_i_pregs_45 : _GEN_1964; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1966 = 7'h2e == io_i_rename_table_15 ? io_i_pregs_46 : _GEN_1965; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1967 = 7'h2f == io_i_rename_table_15 ? io_i_pregs_47 : _GEN_1966; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1968 = 7'h30 == io_i_rename_table_15 ? io_i_pregs_48 : _GEN_1967; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1969 = 7'h31 == io_i_rename_table_15 ? io_i_pregs_49 : _GEN_1968; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1970 = 7'h32 == io_i_rename_table_15 ? io_i_pregs_50 : _GEN_1969; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1971 = 7'h33 == io_i_rename_table_15 ? io_i_pregs_51 : _GEN_1970; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1972 = 7'h34 == io_i_rename_table_15 ? io_i_pregs_52 : _GEN_1971; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1973 = 7'h35 == io_i_rename_table_15 ? io_i_pregs_53 : _GEN_1972; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1974 = 7'h36 == io_i_rename_table_15 ? io_i_pregs_54 : _GEN_1973; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1975 = 7'h37 == io_i_rename_table_15 ? io_i_pregs_55 : _GEN_1974; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1976 = 7'h38 == io_i_rename_table_15 ? io_i_pregs_56 : _GEN_1975; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1977 = 7'h39 == io_i_rename_table_15 ? io_i_pregs_57 : _GEN_1976; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1978 = 7'h3a == io_i_rename_table_15 ? io_i_pregs_58 : _GEN_1977; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1979 = 7'h3b == io_i_rename_table_15 ? io_i_pregs_59 : _GEN_1978; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1980 = 7'h3c == io_i_rename_table_15 ? io_i_pregs_60 : _GEN_1979; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1981 = 7'h3d == io_i_rename_table_15 ? io_i_pregs_61 : _GEN_1980; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1982 = 7'h3e == io_i_rename_table_15 ? io_i_pregs_62 : _GEN_1981; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1983 = 7'h3f == io_i_rename_table_15 ? io_i_pregs_63 : _GEN_1982; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1984 = 7'h40 == io_i_rename_table_15 ? io_i_pregs_64 : _GEN_1983; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1985 = 7'h41 == io_i_rename_table_15 ? io_i_pregs_65 : _GEN_1984; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1986 = 7'h42 == io_i_rename_table_15 ? io_i_pregs_66 : _GEN_1985; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1987 = 7'h43 == io_i_rename_table_15 ? io_i_pregs_67 : _GEN_1986; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1988 = 7'h44 == io_i_rename_table_15 ? io_i_pregs_68 : _GEN_1987; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1989 = 7'h45 == io_i_rename_table_15 ? io_i_pregs_69 : _GEN_1988; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1990 = 7'h46 == io_i_rename_table_15 ? io_i_pregs_70 : _GEN_1989; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1991 = 7'h47 == io_i_rename_table_15 ? io_i_pregs_71 : _GEN_1990; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1992 = 7'h48 == io_i_rename_table_15 ? io_i_pregs_72 : _GEN_1991; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1993 = 7'h49 == io_i_rename_table_15 ? io_i_pregs_73 : _GEN_1992; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1994 = 7'h4a == io_i_rename_table_15 ? io_i_pregs_74 : _GEN_1993; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1995 = 7'h4b == io_i_rename_table_15 ? io_i_pregs_75 : _GEN_1994; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1996 = 7'h4c == io_i_rename_table_15 ? io_i_pregs_76 : _GEN_1995; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1997 = 7'h4d == io_i_rename_table_15 ? io_i_pregs_77 : _GEN_1996; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1998 = 7'h4e == io_i_rename_table_15 ? io_i_pregs_78 : _GEN_1997; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_1999 = 7'h4f == io_i_rename_table_15 ? io_i_pregs_79 : _GEN_1998; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2000 = 7'h50 == io_i_rename_table_15 ? io_i_pregs_80 : _GEN_1999; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2001 = 7'h51 == io_i_rename_table_15 ? io_i_pregs_81 : _GEN_2000; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2002 = 7'h52 == io_i_rename_table_15 ? io_i_pregs_82 : _GEN_2001; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2003 = 7'h53 == io_i_rename_table_15 ? io_i_pregs_83 : _GEN_2002; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2004 = 7'h54 == io_i_rename_table_15 ? io_i_pregs_84 : _GEN_2003; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2005 = 7'h55 == io_i_rename_table_15 ? io_i_pregs_85 : _GEN_2004; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2006 = 7'h56 == io_i_rename_table_15 ? io_i_pregs_86 : _GEN_2005; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2007 = 7'h57 == io_i_rename_table_15 ? io_i_pregs_87 : _GEN_2006; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2008 = 7'h58 == io_i_rename_table_15 ? io_i_pregs_88 : _GEN_2007; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2009 = 7'h59 == io_i_rename_table_15 ? io_i_pregs_89 : _GEN_2008; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2010 = 7'h5a == io_i_rename_table_15 ? io_i_pregs_90 : _GEN_2009; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2011 = 7'h5b == io_i_rename_table_15 ? io_i_pregs_91 : _GEN_2010; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2012 = 7'h5c == io_i_rename_table_15 ? io_i_pregs_92 : _GEN_2011; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2013 = 7'h5d == io_i_rename_table_15 ? io_i_pregs_93 : _GEN_2012; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2014 = 7'h5e == io_i_rename_table_15 ? io_i_pregs_94 : _GEN_2013; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2015 = 7'h5f == io_i_rename_table_15 ? io_i_pregs_95 : _GEN_2014; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2016 = 7'h60 == io_i_rename_table_15 ? io_i_pregs_96 : _GEN_2015; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2017 = 7'h61 == io_i_rename_table_15 ? io_i_pregs_97 : _GEN_2016; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2018 = 7'h62 == io_i_rename_table_15 ? io_i_pregs_98 : _GEN_2017; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2019 = 7'h63 == io_i_rename_table_15 ? io_i_pregs_99 : _GEN_2018; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2020 = 7'h64 == io_i_rename_table_15 ? io_i_pregs_100 : _GEN_2019; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2021 = 7'h65 == io_i_rename_table_15 ? io_i_pregs_101 : _GEN_2020; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2022 = 7'h66 == io_i_rename_table_15 ? io_i_pregs_102 : _GEN_2021; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2023 = 7'h67 == io_i_rename_table_15 ? io_i_pregs_103 : _GEN_2022; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2024 = 7'h68 == io_i_rename_table_15 ? io_i_pregs_104 : _GEN_2023; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2025 = 7'h69 == io_i_rename_table_15 ? io_i_pregs_105 : _GEN_2024; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2026 = 7'h6a == io_i_rename_table_15 ? io_i_pregs_106 : _GEN_2025; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2027 = 7'h6b == io_i_rename_table_15 ? io_i_pregs_107 : _GEN_2026; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2028 = 7'h6c == io_i_rename_table_15 ? io_i_pregs_108 : _GEN_2027; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2029 = 7'h6d == io_i_rename_table_15 ? io_i_pregs_109 : _GEN_2028; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2030 = 7'h6e == io_i_rename_table_15 ? io_i_pregs_110 : _GEN_2029; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2031 = 7'h6f == io_i_rename_table_15 ? io_i_pregs_111 : _GEN_2030; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2032 = 7'h70 == io_i_rename_table_15 ? io_i_pregs_112 : _GEN_2031; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2033 = 7'h71 == io_i_rename_table_15 ? io_i_pregs_113 : _GEN_2032; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2034 = 7'h72 == io_i_rename_table_15 ? io_i_pregs_114 : _GEN_2033; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2035 = 7'h73 == io_i_rename_table_15 ? io_i_pregs_115 : _GEN_2034; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2036 = 7'h74 == io_i_rename_table_15 ? io_i_pregs_116 : _GEN_2035; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2037 = 7'h75 == io_i_rename_table_15 ? io_i_pregs_117 : _GEN_2036; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2038 = 7'h76 == io_i_rename_table_15 ? io_i_pregs_118 : _GEN_2037; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2039 = 7'h77 == io_i_rename_table_15 ? io_i_pregs_119 : _GEN_2038; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2040 = 7'h78 == io_i_rename_table_15 ? io_i_pregs_120 : _GEN_2039; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2041 = 7'h79 == io_i_rename_table_15 ? io_i_pregs_121 : _GEN_2040; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2042 = 7'h7a == io_i_rename_table_15 ? io_i_pregs_122 : _GEN_2041; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2043 = 7'h7b == io_i_rename_table_15 ? io_i_pregs_123 : _GEN_2042; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2044 = 7'h7c == io_i_rename_table_15 ? io_i_pregs_124 : _GEN_2043; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2045 = 7'h7d == io_i_rename_table_15 ? io_i_pregs_125 : _GEN_2044; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2046 = 7'h7e == io_i_rename_table_15 ? io_i_pregs_126 : _GEN_2045; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2049 = 7'h1 == io_i_rename_table_16 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2050 = 7'h2 == io_i_rename_table_16 ? io_i_pregs_2 : _GEN_2049; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2051 = 7'h3 == io_i_rename_table_16 ? io_i_pregs_3 : _GEN_2050; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2052 = 7'h4 == io_i_rename_table_16 ? io_i_pregs_4 : _GEN_2051; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2053 = 7'h5 == io_i_rename_table_16 ? io_i_pregs_5 : _GEN_2052; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2054 = 7'h6 == io_i_rename_table_16 ? io_i_pregs_6 : _GEN_2053; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2055 = 7'h7 == io_i_rename_table_16 ? io_i_pregs_7 : _GEN_2054; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2056 = 7'h8 == io_i_rename_table_16 ? io_i_pregs_8 : _GEN_2055; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2057 = 7'h9 == io_i_rename_table_16 ? io_i_pregs_9 : _GEN_2056; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2058 = 7'ha == io_i_rename_table_16 ? io_i_pregs_10 : _GEN_2057; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2059 = 7'hb == io_i_rename_table_16 ? io_i_pregs_11 : _GEN_2058; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2060 = 7'hc == io_i_rename_table_16 ? io_i_pregs_12 : _GEN_2059; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2061 = 7'hd == io_i_rename_table_16 ? io_i_pregs_13 : _GEN_2060; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2062 = 7'he == io_i_rename_table_16 ? io_i_pregs_14 : _GEN_2061; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2063 = 7'hf == io_i_rename_table_16 ? io_i_pregs_15 : _GEN_2062; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2064 = 7'h10 == io_i_rename_table_16 ? io_i_pregs_16 : _GEN_2063; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2065 = 7'h11 == io_i_rename_table_16 ? io_i_pregs_17 : _GEN_2064; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2066 = 7'h12 == io_i_rename_table_16 ? io_i_pregs_18 : _GEN_2065; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2067 = 7'h13 == io_i_rename_table_16 ? io_i_pregs_19 : _GEN_2066; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2068 = 7'h14 == io_i_rename_table_16 ? io_i_pregs_20 : _GEN_2067; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2069 = 7'h15 == io_i_rename_table_16 ? io_i_pregs_21 : _GEN_2068; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2070 = 7'h16 == io_i_rename_table_16 ? io_i_pregs_22 : _GEN_2069; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2071 = 7'h17 == io_i_rename_table_16 ? io_i_pregs_23 : _GEN_2070; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2072 = 7'h18 == io_i_rename_table_16 ? io_i_pregs_24 : _GEN_2071; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2073 = 7'h19 == io_i_rename_table_16 ? io_i_pregs_25 : _GEN_2072; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2074 = 7'h1a == io_i_rename_table_16 ? io_i_pregs_26 : _GEN_2073; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2075 = 7'h1b == io_i_rename_table_16 ? io_i_pregs_27 : _GEN_2074; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2076 = 7'h1c == io_i_rename_table_16 ? io_i_pregs_28 : _GEN_2075; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2077 = 7'h1d == io_i_rename_table_16 ? io_i_pregs_29 : _GEN_2076; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2078 = 7'h1e == io_i_rename_table_16 ? io_i_pregs_30 : _GEN_2077; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2079 = 7'h1f == io_i_rename_table_16 ? io_i_pregs_31 : _GEN_2078; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2080 = 7'h20 == io_i_rename_table_16 ? io_i_pregs_32 : _GEN_2079; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2081 = 7'h21 == io_i_rename_table_16 ? io_i_pregs_33 : _GEN_2080; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2082 = 7'h22 == io_i_rename_table_16 ? io_i_pregs_34 : _GEN_2081; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2083 = 7'h23 == io_i_rename_table_16 ? io_i_pregs_35 : _GEN_2082; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2084 = 7'h24 == io_i_rename_table_16 ? io_i_pregs_36 : _GEN_2083; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2085 = 7'h25 == io_i_rename_table_16 ? io_i_pregs_37 : _GEN_2084; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2086 = 7'h26 == io_i_rename_table_16 ? io_i_pregs_38 : _GEN_2085; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2087 = 7'h27 == io_i_rename_table_16 ? io_i_pregs_39 : _GEN_2086; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2088 = 7'h28 == io_i_rename_table_16 ? io_i_pregs_40 : _GEN_2087; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2089 = 7'h29 == io_i_rename_table_16 ? io_i_pregs_41 : _GEN_2088; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2090 = 7'h2a == io_i_rename_table_16 ? io_i_pregs_42 : _GEN_2089; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2091 = 7'h2b == io_i_rename_table_16 ? io_i_pregs_43 : _GEN_2090; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2092 = 7'h2c == io_i_rename_table_16 ? io_i_pregs_44 : _GEN_2091; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2093 = 7'h2d == io_i_rename_table_16 ? io_i_pregs_45 : _GEN_2092; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2094 = 7'h2e == io_i_rename_table_16 ? io_i_pregs_46 : _GEN_2093; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2095 = 7'h2f == io_i_rename_table_16 ? io_i_pregs_47 : _GEN_2094; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2096 = 7'h30 == io_i_rename_table_16 ? io_i_pregs_48 : _GEN_2095; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2097 = 7'h31 == io_i_rename_table_16 ? io_i_pregs_49 : _GEN_2096; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2098 = 7'h32 == io_i_rename_table_16 ? io_i_pregs_50 : _GEN_2097; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2099 = 7'h33 == io_i_rename_table_16 ? io_i_pregs_51 : _GEN_2098; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2100 = 7'h34 == io_i_rename_table_16 ? io_i_pregs_52 : _GEN_2099; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2101 = 7'h35 == io_i_rename_table_16 ? io_i_pregs_53 : _GEN_2100; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2102 = 7'h36 == io_i_rename_table_16 ? io_i_pregs_54 : _GEN_2101; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2103 = 7'h37 == io_i_rename_table_16 ? io_i_pregs_55 : _GEN_2102; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2104 = 7'h38 == io_i_rename_table_16 ? io_i_pregs_56 : _GEN_2103; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2105 = 7'h39 == io_i_rename_table_16 ? io_i_pregs_57 : _GEN_2104; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2106 = 7'h3a == io_i_rename_table_16 ? io_i_pregs_58 : _GEN_2105; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2107 = 7'h3b == io_i_rename_table_16 ? io_i_pregs_59 : _GEN_2106; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2108 = 7'h3c == io_i_rename_table_16 ? io_i_pregs_60 : _GEN_2107; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2109 = 7'h3d == io_i_rename_table_16 ? io_i_pregs_61 : _GEN_2108; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2110 = 7'h3e == io_i_rename_table_16 ? io_i_pregs_62 : _GEN_2109; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2111 = 7'h3f == io_i_rename_table_16 ? io_i_pregs_63 : _GEN_2110; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2112 = 7'h40 == io_i_rename_table_16 ? io_i_pregs_64 : _GEN_2111; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2113 = 7'h41 == io_i_rename_table_16 ? io_i_pregs_65 : _GEN_2112; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2114 = 7'h42 == io_i_rename_table_16 ? io_i_pregs_66 : _GEN_2113; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2115 = 7'h43 == io_i_rename_table_16 ? io_i_pregs_67 : _GEN_2114; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2116 = 7'h44 == io_i_rename_table_16 ? io_i_pregs_68 : _GEN_2115; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2117 = 7'h45 == io_i_rename_table_16 ? io_i_pregs_69 : _GEN_2116; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2118 = 7'h46 == io_i_rename_table_16 ? io_i_pregs_70 : _GEN_2117; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2119 = 7'h47 == io_i_rename_table_16 ? io_i_pregs_71 : _GEN_2118; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2120 = 7'h48 == io_i_rename_table_16 ? io_i_pregs_72 : _GEN_2119; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2121 = 7'h49 == io_i_rename_table_16 ? io_i_pregs_73 : _GEN_2120; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2122 = 7'h4a == io_i_rename_table_16 ? io_i_pregs_74 : _GEN_2121; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2123 = 7'h4b == io_i_rename_table_16 ? io_i_pregs_75 : _GEN_2122; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2124 = 7'h4c == io_i_rename_table_16 ? io_i_pregs_76 : _GEN_2123; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2125 = 7'h4d == io_i_rename_table_16 ? io_i_pregs_77 : _GEN_2124; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2126 = 7'h4e == io_i_rename_table_16 ? io_i_pregs_78 : _GEN_2125; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2127 = 7'h4f == io_i_rename_table_16 ? io_i_pregs_79 : _GEN_2126; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2128 = 7'h50 == io_i_rename_table_16 ? io_i_pregs_80 : _GEN_2127; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2129 = 7'h51 == io_i_rename_table_16 ? io_i_pregs_81 : _GEN_2128; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2130 = 7'h52 == io_i_rename_table_16 ? io_i_pregs_82 : _GEN_2129; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2131 = 7'h53 == io_i_rename_table_16 ? io_i_pregs_83 : _GEN_2130; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2132 = 7'h54 == io_i_rename_table_16 ? io_i_pregs_84 : _GEN_2131; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2133 = 7'h55 == io_i_rename_table_16 ? io_i_pregs_85 : _GEN_2132; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2134 = 7'h56 == io_i_rename_table_16 ? io_i_pregs_86 : _GEN_2133; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2135 = 7'h57 == io_i_rename_table_16 ? io_i_pregs_87 : _GEN_2134; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2136 = 7'h58 == io_i_rename_table_16 ? io_i_pregs_88 : _GEN_2135; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2137 = 7'h59 == io_i_rename_table_16 ? io_i_pregs_89 : _GEN_2136; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2138 = 7'h5a == io_i_rename_table_16 ? io_i_pregs_90 : _GEN_2137; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2139 = 7'h5b == io_i_rename_table_16 ? io_i_pregs_91 : _GEN_2138; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2140 = 7'h5c == io_i_rename_table_16 ? io_i_pregs_92 : _GEN_2139; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2141 = 7'h5d == io_i_rename_table_16 ? io_i_pregs_93 : _GEN_2140; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2142 = 7'h5e == io_i_rename_table_16 ? io_i_pregs_94 : _GEN_2141; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2143 = 7'h5f == io_i_rename_table_16 ? io_i_pregs_95 : _GEN_2142; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2144 = 7'h60 == io_i_rename_table_16 ? io_i_pregs_96 : _GEN_2143; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2145 = 7'h61 == io_i_rename_table_16 ? io_i_pregs_97 : _GEN_2144; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2146 = 7'h62 == io_i_rename_table_16 ? io_i_pregs_98 : _GEN_2145; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2147 = 7'h63 == io_i_rename_table_16 ? io_i_pregs_99 : _GEN_2146; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2148 = 7'h64 == io_i_rename_table_16 ? io_i_pregs_100 : _GEN_2147; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2149 = 7'h65 == io_i_rename_table_16 ? io_i_pregs_101 : _GEN_2148; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2150 = 7'h66 == io_i_rename_table_16 ? io_i_pregs_102 : _GEN_2149; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2151 = 7'h67 == io_i_rename_table_16 ? io_i_pregs_103 : _GEN_2150; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2152 = 7'h68 == io_i_rename_table_16 ? io_i_pregs_104 : _GEN_2151; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2153 = 7'h69 == io_i_rename_table_16 ? io_i_pregs_105 : _GEN_2152; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2154 = 7'h6a == io_i_rename_table_16 ? io_i_pregs_106 : _GEN_2153; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2155 = 7'h6b == io_i_rename_table_16 ? io_i_pregs_107 : _GEN_2154; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2156 = 7'h6c == io_i_rename_table_16 ? io_i_pregs_108 : _GEN_2155; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2157 = 7'h6d == io_i_rename_table_16 ? io_i_pregs_109 : _GEN_2156; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2158 = 7'h6e == io_i_rename_table_16 ? io_i_pregs_110 : _GEN_2157; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2159 = 7'h6f == io_i_rename_table_16 ? io_i_pregs_111 : _GEN_2158; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2160 = 7'h70 == io_i_rename_table_16 ? io_i_pregs_112 : _GEN_2159; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2161 = 7'h71 == io_i_rename_table_16 ? io_i_pregs_113 : _GEN_2160; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2162 = 7'h72 == io_i_rename_table_16 ? io_i_pregs_114 : _GEN_2161; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2163 = 7'h73 == io_i_rename_table_16 ? io_i_pregs_115 : _GEN_2162; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2164 = 7'h74 == io_i_rename_table_16 ? io_i_pregs_116 : _GEN_2163; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2165 = 7'h75 == io_i_rename_table_16 ? io_i_pregs_117 : _GEN_2164; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2166 = 7'h76 == io_i_rename_table_16 ? io_i_pregs_118 : _GEN_2165; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2167 = 7'h77 == io_i_rename_table_16 ? io_i_pregs_119 : _GEN_2166; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2168 = 7'h78 == io_i_rename_table_16 ? io_i_pregs_120 : _GEN_2167; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2169 = 7'h79 == io_i_rename_table_16 ? io_i_pregs_121 : _GEN_2168; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2170 = 7'h7a == io_i_rename_table_16 ? io_i_pregs_122 : _GEN_2169; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2171 = 7'h7b == io_i_rename_table_16 ? io_i_pregs_123 : _GEN_2170; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2172 = 7'h7c == io_i_rename_table_16 ? io_i_pregs_124 : _GEN_2171; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2173 = 7'h7d == io_i_rename_table_16 ? io_i_pregs_125 : _GEN_2172; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2174 = 7'h7e == io_i_rename_table_16 ? io_i_pregs_126 : _GEN_2173; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2177 = 7'h1 == io_i_rename_table_17 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2178 = 7'h2 == io_i_rename_table_17 ? io_i_pregs_2 : _GEN_2177; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2179 = 7'h3 == io_i_rename_table_17 ? io_i_pregs_3 : _GEN_2178; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2180 = 7'h4 == io_i_rename_table_17 ? io_i_pregs_4 : _GEN_2179; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2181 = 7'h5 == io_i_rename_table_17 ? io_i_pregs_5 : _GEN_2180; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2182 = 7'h6 == io_i_rename_table_17 ? io_i_pregs_6 : _GEN_2181; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2183 = 7'h7 == io_i_rename_table_17 ? io_i_pregs_7 : _GEN_2182; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2184 = 7'h8 == io_i_rename_table_17 ? io_i_pregs_8 : _GEN_2183; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2185 = 7'h9 == io_i_rename_table_17 ? io_i_pregs_9 : _GEN_2184; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2186 = 7'ha == io_i_rename_table_17 ? io_i_pregs_10 : _GEN_2185; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2187 = 7'hb == io_i_rename_table_17 ? io_i_pregs_11 : _GEN_2186; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2188 = 7'hc == io_i_rename_table_17 ? io_i_pregs_12 : _GEN_2187; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2189 = 7'hd == io_i_rename_table_17 ? io_i_pregs_13 : _GEN_2188; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2190 = 7'he == io_i_rename_table_17 ? io_i_pregs_14 : _GEN_2189; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2191 = 7'hf == io_i_rename_table_17 ? io_i_pregs_15 : _GEN_2190; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2192 = 7'h10 == io_i_rename_table_17 ? io_i_pregs_16 : _GEN_2191; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2193 = 7'h11 == io_i_rename_table_17 ? io_i_pregs_17 : _GEN_2192; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2194 = 7'h12 == io_i_rename_table_17 ? io_i_pregs_18 : _GEN_2193; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2195 = 7'h13 == io_i_rename_table_17 ? io_i_pregs_19 : _GEN_2194; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2196 = 7'h14 == io_i_rename_table_17 ? io_i_pregs_20 : _GEN_2195; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2197 = 7'h15 == io_i_rename_table_17 ? io_i_pregs_21 : _GEN_2196; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2198 = 7'h16 == io_i_rename_table_17 ? io_i_pregs_22 : _GEN_2197; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2199 = 7'h17 == io_i_rename_table_17 ? io_i_pregs_23 : _GEN_2198; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2200 = 7'h18 == io_i_rename_table_17 ? io_i_pregs_24 : _GEN_2199; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2201 = 7'h19 == io_i_rename_table_17 ? io_i_pregs_25 : _GEN_2200; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2202 = 7'h1a == io_i_rename_table_17 ? io_i_pregs_26 : _GEN_2201; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2203 = 7'h1b == io_i_rename_table_17 ? io_i_pregs_27 : _GEN_2202; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2204 = 7'h1c == io_i_rename_table_17 ? io_i_pregs_28 : _GEN_2203; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2205 = 7'h1d == io_i_rename_table_17 ? io_i_pregs_29 : _GEN_2204; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2206 = 7'h1e == io_i_rename_table_17 ? io_i_pregs_30 : _GEN_2205; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2207 = 7'h1f == io_i_rename_table_17 ? io_i_pregs_31 : _GEN_2206; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2208 = 7'h20 == io_i_rename_table_17 ? io_i_pregs_32 : _GEN_2207; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2209 = 7'h21 == io_i_rename_table_17 ? io_i_pregs_33 : _GEN_2208; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2210 = 7'h22 == io_i_rename_table_17 ? io_i_pregs_34 : _GEN_2209; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2211 = 7'h23 == io_i_rename_table_17 ? io_i_pregs_35 : _GEN_2210; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2212 = 7'h24 == io_i_rename_table_17 ? io_i_pregs_36 : _GEN_2211; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2213 = 7'h25 == io_i_rename_table_17 ? io_i_pregs_37 : _GEN_2212; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2214 = 7'h26 == io_i_rename_table_17 ? io_i_pregs_38 : _GEN_2213; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2215 = 7'h27 == io_i_rename_table_17 ? io_i_pregs_39 : _GEN_2214; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2216 = 7'h28 == io_i_rename_table_17 ? io_i_pregs_40 : _GEN_2215; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2217 = 7'h29 == io_i_rename_table_17 ? io_i_pregs_41 : _GEN_2216; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2218 = 7'h2a == io_i_rename_table_17 ? io_i_pregs_42 : _GEN_2217; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2219 = 7'h2b == io_i_rename_table_17 ? io_i_pregs_43 : _GEN_2218; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2220 = 7'h2c == io_i_rename_table_17 ? io_i_pregs_44 : _GEN_2219; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2221 = 7'h2d == io_i_rename_table_17 ? io_i_pregs_45 : _GEN_2220; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2222 = 7'h2e == io_i_rename_table_17 ? io_i_pregs_46 : _GEN_2221; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2223 = 7'h2f == io_i_rename_table_17 ? io_i_pregs_47 : _GEN_2222; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2224 = 7'h30 == io_i_rename_table_17 ? io_i_pregs_48 : _GEN_2223; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2225 = 7'h31 == io_i_rename_table_17 ? io_i_pregs_49 : _GEN_2224; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2226 = 7'h32 == io_i_rename_table_17 ? io_i_pregs_50 : _GEN_2225; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2227 = 7'h33 == io_i_rename_table_17 ? io_i_pregs_51 : _GEN_2226; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2228 = 7'h34 == io_i_rename_table_17 ? io_i_pregs_52 : _GEN_2227; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2229 = 7'h35 == io_i_rename_table_17 ? io_i_pregs_53 : _GEN_2228; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2230 = 7'h36 == io_i_rename_table_17 ? io_i_pregs_54 : _GEN_2229; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2231 = 7'h37 == io_i_rename_table_17 ? io_i_pregs_55 : _GEN_2230; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2232 = 7'h38 == io_i_rename_table_17 ? io_i_pregs_56 : _GEN_2231; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2233 = 7'h39 == io_i_rename_table_17 ? io_i_pregs_57 : _GEN_2232; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2234 = 7'h3a == io_i_rename_table_17 ? io_i_pregs_58 : _GEN_2233; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2235 = 7'h3b == io_i_rename_table_17 ? io_i_pregs_59 : _GEN_2234; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2236 = 7'h3c == io_i_rename_table_17 ? io_i_pregs_60 : _GEN_2235; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2237 = 7'h3d == io_i_rename_table_17 ? io_i_pregs_61 : _GEN_2236; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2238 = 7'h3e == io_i_rename_table_17 ? io_i_pregs_62 : _GEN_2237; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2239 = 7'h3f == io_i_rename_table_17 ? io_i_pregs_63 : _GEN_2238; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2240 = 7'h40 == io_i_rename_table_17 ? io_i_pregs_64 : _GEN_2239; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2241 = 7'h41 == io_i_rename_table_17 ? io_i_pregs_65 : _GEN_2240; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2242 = 7'h42 == io_i_rename_table_17 ? io_i_pregs_66 : _GEN_2241; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2243 = 7'h43 == io_i_rename_table_17 ? io_i_pregs_67 : _GEN_2242; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2244 = 7'h44 == io_i_rename_table_17 ? io_i_pregs_68 : _GEN_2243; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2245 = 7'h45 == io_i_rename_table_17 ? io_i_pregs_69 : _GEN_2244; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2246 = 7'h46 == io_i_rename_table_17 ? io_i_pregs_70 : _GEN_2245; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2247 = 7'h47 == io_i_rename_table_17 ? io_i_pregs_71 : _GEN_2246; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2248 = 7'h48 == io_i_rename_table_17 ? io_i_pregs_72 : _GEN_2247; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2249 = 7'h49 == io_i_rename_table_17 ? io_i_pregs_73 : _GEN_2248; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2250 = 7'h4a == io_i_rename_table_17 ? io_i_pregs_74 : _GEN_2249; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2251 = 7'h4b == io_i_rename_table_17 ? io_i_pregs_75 : _GEN_2250; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2252 = 7'h4c == io_i_rename_table_17 ? io_i_pregs_76 : _GEN_2251; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2253 = 7'h4d == io_i_rename_table_17 ? io_i_pregs_77 : _GEN_2252; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2254 = 7'h4e == io_i_rename_table_17 ? io_i_pregs_78 : _GEN_2253; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2255 = 7'h4f == io_i_rename_table_17 ? io_i_pregs_79 : _GEN_2254; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2256 = 7'h50 == io_i_rename_table_17 ? io_i_pregs_80 : _GEN_2255; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2257 = 7'h51 == io_i_rename_table_17 ? io_i_pregs_81 : _GEN_2256; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2258 = 7'h52 == io_i_rename_table_17 ? io_i_pregs_82 : _GEN_2257; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2259 = 7'h53 == io_i_rename_table_17 ? io_i_pregs_83 : _GEN_2258; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2260 = 7'h54 == io_i_rename_table_17 ? io_i_pregs_84 : _GEN_2259; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2261 = 7'h55 == io_i_rename_table_17 ? io_i_pregs_85 : _GEN_2260; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2262 = 7'h56 == io_i_rename_table_17 ? io_i_pregs_86 : _GEN_2261; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2263 = 7'h57 == io_i_rename_table_17 ? io_i_pregs_87 : _GEN_2262; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2264 = 7'h58 == io_i_rename_table_17 ? io_i_pregs_88 : _GEN_2263; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2265 = 7'h59 == io_i_rename_table_17 ? io_i_pregs_89 : _GEN_2264; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2266 = 7'h5a == io_i_rename_table_17 ? io_i_pregs_90 : _GEN_2265; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2267 = 7'h5b == io_i_rename_table_17 ? io_i_pregs_91 : _GEN_2266; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2268 = 7'h5c == io_i_rename_table_17 ? io_i_pregs_92 : _GEN_2267; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2269 = 7'h5d == io_i_rename_table_17 ? io_i_pregs_93 : _GEN_2268; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2270 = 7'h5e == io_i_rename_table_17 ? io_i_pregs_94 : _GEN_2269; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2271 = 7'h5f == io_i_rename_table_17 ? io_i_pregs_95 : _GEN_2270; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2272 = 7'h60 == io_i_rename_table_17 ? io_i_pregs_96 : _GEN_2271; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2273 = 7'h61 == io_i_rename_table_17 ? io_i_pregs_97 : _GEN_2272; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2274 = 7'h62 == io_i_rename_table_17 ? io_i_pregs_98 : _GEN_2273; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2275 = 7'h63 == io_i_rename_table_17 ? io_i_pregs_99 : _GEN_2274; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2276 = 7'h64 == io_i_rename_table_17 ? io_i_pregs_100 : _GEN_2275; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2277 = 7'h65 == io_i_rename_table_17 ? io_i_pregs_101 : _GEN_2276; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2278 = 7'h66 == io_i_rename_table_17 ? io_i_pregs_102 : _GEN_2277; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2279 = 7'h67 == io_i_rename_table_17 ? io_i_pregs_103 : _GEN_2278; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2280 = 7'h68 == io_i_rename_table_17 ? io_i_pregs_104 : _GEN_2279; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2281 = 7'h69 == io_i_rename_table_17 ? io_i_pregs_105 : _GEN_2280; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2282 = 7'h6a == io_i_rename_table_17 ? io_i_pregs_106 : _GEN_2281; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2283 = 7'h6b == io_i_rename_table_17 ? io_i_pregs_107 : _GEN_2282; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2284 = 7'h6c == io_i_rename_table_17 ? io_i_pregs_108 : _GEN_2283; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2285 = 7'h6d == io_i_rename_table_17 ? io_i_pregs_109 : _GEN_2284; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2286 = 7'h6e == io_i_rename_table_17 ? io_i_pregs_110 : _GEN_2285; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2287 = 7'h6f == io_i_rename_table_17 ? io_i_pregs_111 : _GEN_2286; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2288 = 7'h70 == io_i_rename_table_17 ? io_i_pregs_112 : _GEN_2287; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2289 = 7'h71 == io_i_rename_table_17 ? io_i_pregs_113 : _GEN_2288; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2290 = 7'h72 == io_i_rename_table_17 ? io_i_pregs_114 : _GEN_2289; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2291 = 7'h73 == io_i_rename_table_17 ? io_i_pregs_115 : _GEN_2290; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2292 = 7'h74 == io_i_rename_table_17 ? io_i_pregs_116 : _GEN_2291; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2293 = 7'h75 == io_i_rename_table_17 ? io_i_pregs_117 : _GEN_2292; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2294 = 7'h76 == io_i_rename_table_17 ? io_i_pregs_118 : _GEN_2293; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2295 = 7'h77 == io_i_rename_table_17 ? io_i_pregs_119 : _GEN_2294; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2296 = 7'h78 == io_i_rename_table_17 ? io_i_pregs_120 : _GEN_2295; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2297 = 7'h79 == io_i_rename_table_17 ? io_i_pregs_121 : _GEN_2296; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2298 = 7'h7a == io_i_rename_table_17 ? io_i_pregs_122 : _GEN_2297; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2299 = 7'h7b == io_i_rename_table_17 ? io_i_pregs_123 : _GEN_2298; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2300 = 7'h7c == io_i_rename_table_17 ? io_i_pregs_124 : _GEN_2299; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2301 = 7'h7d == io_i_rename_table_17 ? io_i_pregs_125 : _GEN_2300; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2302 = 7'h7e == io_i_rename_table_17 ? io_i_pregs_126 : _GEN_2301; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2305 = 7'h1 == io_i_rename_table_18 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2306 = 7'h2 == io_i_rename_table_18 ? io_i_pregs_2 : _GEN_2305; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2307 = 7'h3 == io_i_rename_table_18 ? io_i_pregs_3 : _GEN_2306; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2308 = 7'h4 == io_i_rename_table_18 ? io_i_pregs_4 : _GEN_2307; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2309 = 7'h5 == io_i_rename_table_18 ? io_i_pregs_5 : _GEN_2308; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2310 = 7'h6 == io_i_rename_table_18 ? io_i_pregs_6 : _GEN_2309; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2311 = 7'h7 == io_i_rename_table_18 ? io_i_pregs_7 : _GEN_2310; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2312 = 7'h8 == io_i_rename_table_18 ? io_i_pregs_8 : _GEN_2311; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2313 = 7'h9 == io_i_rename_table_18 ? io_i_pregs_9 : _GEN_2312; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2314 = 7'ha == io_i_rename_table_18 ? io_i_pregs_10 : _GEN_2313; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2315 = 7'hb == io_i_rename_table_18 ? io_i_pregs_11 : _GEN_2314; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2316 = 7'hc == io_i_rename_table_18 ? io_i_pregs_12 : _GEN_2315; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2317 = 7'hd == io_i_rename_table_18 ? io_i_pregs_13 : _GEN_2316; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2318 = 7'he == io_i_rename_table_18 ? io_i_pregs_14 : _GEN_2317; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2319 = 7'hf == io_i_rename_table_18 ? io_i_pregs_15 : _GEN_2318; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2320 = 7'h10 == io_i_rename_table_18 ? io_i_pregs_16 : _GEN_2319; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2321 = 7'h11 == io_i_rename_table_18 ? io_i_pregs_17 : _GEN_2320; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2322 = 7'h12 == io_i_rename_table_18 ? io_i_pregs_18 : _GEN_2321; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2323 = 7'h13 == io_i_rename_table_18 ? io_i_pregs_19 : _GEN_2322; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2324 = 7'h14 == io_i_rename_table_18 ? io_i_pregs_20 : _GEN_2323; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2325 = 7'h15 == io_i_rename_table_18 ? io_i_pregs_21 : _GEN_2324; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2326 = 7'h16 == io_i_rename_table_18 ? io_i_pregs_22 : _GEN_2325; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2327 = 7'h17 == io_i_rename_table_18 ? io_i_pregs_23 : _GEN_2326; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2328 = 7'h18 == io_i_rename_table_18 ? io_i_pregs_24 : _GEN_2327; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2329 = 7'h19 == io_i_rename_table_18 ? io_i_pregs_25 : _GEN_2328; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2330 = 7'h1a == io_i_rename_table_18 ? io_i_pregs_26 : _GEN_2329; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2331 = 7'h1b == io_i_rename_table_18 ? io_i_pregs_27 : _GEN_2330; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2332 = 7'h1c == io_i_rename_table_18 ? io_i_pregs_28 : _GEN_2331; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2333 = 7'h1d == io_i_rename_table_18 ? io_i_pregs_29 : _GEN_2332; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2334 = 7'h1e == io_i_rename_table_18 ? io_i_pregs_30 : _GEN_2333; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2335 = 7'h1f == io_i_rename_table_18 ? io_i_pregs_31 : _GEN_2334; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2336 = 7'h20 == io_i_rename_table_18 ? io_i_pregs_32 : _GEN_2335; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2337 = 7'h21 == io_i_rename_table_18 ? io_i_pregs_33 : _GEN_2336; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2338 = 7'h22 == io_i_rename_table_18 ? io_i_pregs_34 : _GEN_2337; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2339 = 7'h23 == io_i_rename_table_18 ? io_i_pregs_35 : _GEN_2338; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2340 = 7'h24 == io_i_rename_table_18 ? io_i_pregs_36 : _GEN_2339; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2341 = 7'h25 == io_i_rename_table_18 ? io_i_pregs_37 : _GEN_2340; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2342 = 7'h26 == io_i_rename_table_18 ? io_i_pregs_38 : _GEN_2341; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2343 = 7'h27 == io_i_rename_table_18 ? io_i_pregs_39 : _GEN_2342; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2344 = 7'h28 == io_i_rename_table_18 ? io_i_pregs_40 : _GEN_2343; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2345 = 7'h29 == io_i_rename_table_18 ? io_i_pregs_41 : _GEN_2344; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2346 = 7'h2a == io_i_rename_table_18 ? io_i_pregs_42 : _GEN_2345; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2347 = 7'h2b == io_i_rename_table_18 ? io_i_pregs_43 : _GEN_2346; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2348 = 7'h2c == io_i_rename_table_18 ? io_i_pregs_44 : _GEN_2347; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2349 = 7'h2d == io_i_rename_table_18 ? io_i_pregs_45 : _GEN_2348; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2350 = 7'h2e == io_i_rename_table_18 ? io_i_pregs_46 : _GEN_2349; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2351 = 7'h2f == io_i_rename_table_18 ? io_i_pregs_47 : _GEN_2350; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2352 = 7'h30 == io_i_rename_table_18 ? io_i_pregs_48 : _GEN_2351; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2353 = 7'h31 == io_i_rename_table_18 ? io_i_pregs_49 : _GEN_2352; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2354 = 7'h32 == io_i_rename_table_18 ? io_i_pregs_50 : _GEN_2353; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2355 = 7'h33 == io_i_rename_table_18 ? io_i_pregs_51 : _GEN_2354; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2356 = 7'h34 == io_i_rename_table_18 ? io_i_pregs_52 : _GEN_2355; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2357 = 7'h35 == io_i_rename_table_18 ? io_i_pregs_53 : _GEN_2356; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2358 = 7'h36 == io_i_rename_table_18 ? io_i_pregs_54 : _GEN_2357; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2359 = 7'h37 == io_i_rename_table_18 ? io_i_pregs_55 : _GEN_2358; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2360 = 7'h38 == io_i_rename_table_18 ? io_i_pregs_56 : _GEN_2359; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2361 = 7'h39 == io_i_rename_table_18 ? io_i_pregs_57 : _GEN_2360; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2362 = 7'h3a == io_i_rename_table_18 ? io_i_pregs_58 : _GEN_2361; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2363 = 7'h3b == io_i_rename_table_18 ? io_i_pregs_59 : _GEN_2362; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2364 = 7'h3c == io_i_rename_table_18 ? io_i_pregs_60 : _GEN_2363; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2365 = 7'h3d == io_i_rename_table_18 ? io_i_pregs_61 : _GEN_2364; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2366 = 7'h3e == io_i_rename_table_18 ? io_i_pregs_62 : _GEN_2365; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2367 = 7'h3f == io_i_rename_table_18 ? io_i_pregs_63 : _GEN_2366; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2368 = 7'h40 == io_i_rename_table_18 ? io_i_pregs_64 : _GEN_2367; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2369 = 7'h41 == io_i_rename_table_18 ? io_i_pregs_65 : _GEN_2368; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2370 = 7'h42 == io_i_rename_table_18 ? io_i_pregs_66 : _GEN_2369; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2371 = 7'h43 == io_i_rename_table_18 ? io_i_pregs_67 : _GEN_2370; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2372 = 7'h44 == io_i_rename_table_18 ? io_i_pregs_68 : _GEN_2371; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2373 = 7'h45 == io_i_rename_table_18 ? io_i_pregs_69 : _GEN_2372; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2374 = 7'h46 == io_i_rename_table_18 ? io_i_pregs_70 : _GEN_2373; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2375 = 7'h47 == io_i_rename_table_18 ? io_i_pregs_71 : _GEN_2374; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2376 = 7'h48 == io_i_rename_table_18 ? io_i_pregs_72 : _GEN_2375; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2377 = 7'h49 == io_i_rename_table_18 ? io_i_pregs_73 : _GEN_2376; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2378 = 7'h4a == io_i_rename_table_18 ? io_i_pregs_74 : _GEN_2377; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2379 = 7'h4b == io_i_rename_table_18 ? io_i_pregs_75 : _GEN_2378; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2380 = 7'h4c == io_i_rename_table_18 ? io_i_pregs_76 : _GEN_2379; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2381 = 7'h4d == io_i_rename_table_18 ? io_i_pregs_77 : _GEN_2380; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2382 = 7'h4e == io_i_rename_table_18 ? io_i_pregs_78 : _GEN_2381; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2383 = 7'h4f == io_i_rename_table_18 ? io_i_pregs_79 : _GEN_2382; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2384 = 7'h50 == io_i_rename_table_18 ? io_i_pregs_80 : _GEN_2383; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2385 = 7'h51 == io_i_rename_table_18 ? io_i_pregs_81 : _GEN_2384; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2386 = 7'h52 == io_i_rename_table_18 ? io_i_pregs_82 : _GEN_2385; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2387 = 7'h53 == io_i_rename_table_18 ? io_i_pregs_83 : _GEN_2386; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2388 = 7'h54 == io_i_rename_table_18 ? io_i_pregs_84 : _GEN_2387; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2389 = 7'h55 == io_i_rename_table_18 ? io_i_pregs_85 : _GEN_2388; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2390 = 7'h56 == io_i_rename_table_18 ? io_i_pregs_86 : _GEN_2389; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2391 = 7'h57 == io_i_rename_table_18 ? io_i_pregs_87 : _GEN_2390; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2392 = 7'h58 == io_i_rename_table_18 ? io_i_pregs_88 : _GEN_2391; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2393 = 7'h59 == io_i_rename_table_18 ? io_i_pregs_89 : _GEN_2392; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2394 = 7'h5a == io_i_rename_table_18 ? io_i_pregs_90 : _GEN_2393; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2395 = 7'h5b == io_i_rename_table_18 ? io_i_pregs_91 : _GEN_2394; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2396 = 7'h5c == io_i_rename_table_18 ? io_i_pregs_92 : _GEN_2395; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2397 = 7'h5d == io_i_rename_table_18 ? io_i_pregs_93 : _GEN_2396; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2398 = 7'h5e == io_i_rename_table_18 ? io_i_pregs_94 : _GEN_2397; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2399 = 7'h5f == io_i_rename_table_18 ? io_i_pregs_95 : _GEN_2398; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2400 = 7'h60 == io_i_rename_table_18 ? io_i_pregs_96 : _GEN_2399; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2401 = 7'h61 == io_i_rename_table_18 ? io_i_pregs_97 : _GEN_2400; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2402 = 7'h62 == io_i_rename_table_18 ? io_i_pregs_98 : _GEN_2401; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2403 = 7'h63 == io_i_rename_table_18 ? io_i_pregs_99 : _GEN_2402; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2404 = 7'h64 == io_i_rename_table_18 ? io_i_pregs_100 : _GEN_2403; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2405 = 7'h65 == io_i_rename_table_18 ? io_i_pregs_101 : _GEN_2404; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2406 = 7'h66 == io_i_rename_table_18 ? io_i_pregs_102 : _GEN_2405; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2407 = 7'h67 == io_i_rename_table_18 ? io_i_pregs_103 : _GEN_2406; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2408 = 7'h68 == io_i_rename_table_18 ? io_i_pregs_104 : _GEN_2407; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2409 = 7'h69 == io_i_rename_table_18 ? io_i_pregs_105 : _GEN_2408; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2410 = 7'h6a == io_i_rename_table_18 ? io_i_pregs_106 : _GEN_2409; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2411 = 7'h6b == io_i_rename_table_18 ? io_i_pregs_107 : _GEN_2410; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2412 = 7'h6c == io_i_rename_table_18 ? io_i_pregs_108 : _GEN_2411; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2413 = 7'h6d == io_i_rename_table_18 ? io_i_pregs_109 : _GEN_2412; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2414 = 7'h6e == io_i_rename_table_18 ? io_i_pregs_110 : _GEN_2413; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2415 = 7'h6f == io_i_rename_table_18 ? io_i_pregs_111 : _GEN_2414; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2416 = 7'h70 == io_i_rename_table_18 ? io_i_pregs_112 : _GEN_2415; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2417 = 7'h71 == io_i_rename_table_18 ? io_i_pregs_113 : _GEN_2416; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2418 = 7'h72 == io_i_rename_table_18 ? io_i_pregs_114 : _GEN_2417; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2419 = 7'h73 == io_i_rename_table_18 ? io_i_pregs_115 : _GEN_2418; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2420 = 7'h74 == io_i_rename_table_18 ? io_i_pregs_116 : _GEN_2419; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2421 = 7'h75 == io_i_rename_table_18 ? io_i_pregs_117 : _GEN_2420; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2422 = 7'h76 == io_i_rename_table_18 ? io_i_pregs_118 : _GEN_2421; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2423 = 7'h77 == io_i_rename_table_18 ? io_i_pregs_119 : _GEN_2422; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2424 = 7'h78 == io_i_rename_table_18 ? io_i_pregs_120 : _GEN_2423; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2425 = 7'h79 == io_i_rename_table_18 ? io_i_pregs_121 : _GEN_2424; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2426 = 7'h7a == io_i_rename_table_18 ? io_i_pregs_122 : _GEN_2425; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2427 = 7'h7b == io_i_rename_table_18 ? io_i_pregs_123 : _GEN_2426; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2428 = 7'h7c == io_i_rename_table_18 ? io_i_pregs_124 : _GEN_2427; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2429 = 7'h7d == io_i_rename_table_18 ? io_i_pregs_125 : _GEN_2428; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2430 = 7'h7e == io_i_rename_table_18 ? io_i_pregs_126 : _GEN_2429; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2433 = 7'h1 == io_i_rename_table_19 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2434 = 7'h2 == io_i_rename_table_19 ? io_i_pregs_2 : _GEN_2433; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2435 = 7'h3 == io_i_rename_table_19 ? io_i_pregs_3 : _GEN_2434; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2436 = 7'h4 == io_i_rename_table_19 ? io_i_pregs_4 : _GEN_2435; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2437 = 7'h5 == io_i_rename_table_19 ? io_i_pregs_5 : _GEN_2436; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2438 = 7'h6 == io_i_rename_table_19 ? io_i_pregs_6 : _GEN_2437; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2439 = 7'h7 == io_i_rename_table_19 ? io_i_pregs_7 : _GEN_2438; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2440 = 7'h8 == io_i_rename_table_19 ? io_i_pregs_8 : _GEN_2439; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2441 = 7'h9 == io_i_rename_table_19 ? io_i_pregs_9 : _GEN_2440; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2442 = 7'ha == io_i_rename_table_19 ? io_i_pregs_10 : _GEN_2441; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2443 = 7'hb == io_i_rename_table_19 ? io_i_pregs_11 : _GEN_2442; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2444 = 7'hc == io_i_rename_table_19 ? io_i_pregs_12 : _GEN_2443; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2445 = 7'hd == io_i_rename_table_19 ? io_i_pregs_13 : _GEN_2444; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2446 = 7'he == io_i_rename_table_19 ? io_i_pregs_14 : _GEN_2445; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2447 = 7'hf == io_i_rename_table_19 ? io_i_pregs_15 : _GEN_2446; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2448 = 7'h10 == io_i_rename_table_19 ? io_i_pregs_16 : _GEN_2447; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2449 = 7'h11 == io_i_rename_table_19 ? io_i_pregs_17 : _GEN_2448; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2450 = 7'h12 == io_i_rename_table_19 ? io_i_pregs_18 : _GEN_2449; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2451 = 7'h13 == io_i_rename_table_19 ? io_i_pregs_19 : _GEN_2450; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2452 = 7'h14 == io_i_rename_table_19 ? io_i_pregs_20 : _GEN_2451; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2453 = 7'h15 == io_i_rename_table_19 ? io_i_pregs_21 : _GEN_2452; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2454 = 7'h16 == io_i_rename_table_19 ? io_i_pregs_22 : _GEN_2453; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2455 = 7'h17 == io_i_rename_table_19 ? io_i_pregs_23 : _GEN_2454; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2456 = 7'h18 == io_i_rename_table_19 ? io_i_pregs_24 : _GEN_2455; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2457 = 7'h19 == io_i_rename_table_19 ? io_i_pregs_25 : _GEN_2456; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2458 = 7'h1a == io_i_rename_table_19 ? io_i_pregs_26 : _GEN_2457; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2459 = 7'h1b == io_i_rename_table_19 ? io_i_pregs_27 : _GEN_2458; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2460 = 7'h1c == io_i_rename_table_19 ? io_i_pregs_28 : _GEN_2459; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2461 = 7'h1d == io_i_rename_table_19 ? io_i_pregs_29 : _GEN_2460; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2462 = 7'h1e == io_i_rename_table_19 ? io_i_pregs_30 : _GEN_2461; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2463 = 7'h1f == io_i_rename_table_19 ? io_i_pregs_31 : _GEN_2462; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2464 = 7'h20 == io_i_rename_table_19 ? io_i_pregs_32 : _GEN_2463; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2465 = 7'h21 == io_i_rename_table_19 ? io_i_pregs_33 : _GEN_2464; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2466 = 7'h22 == io_i_rename_table_19 ? io_i_pregs_34 : _GEN_2465; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2467 = 7'h23 == io_i_rename_table_19 ? io_i_pregs_35 : _GEN_2466; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2468 = 7'h24 == io_i_rename_table_19 ? io_i_pregs_36 : _GEN_2467; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2469 = 7'h25 == io_i_rename_table_19 ? io_i_pregs_37 : _GEN_2468; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2470 = 7'h26 == io_i_rename_table_19 ? io_i_pregs_38 : _GEN_2469; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2471 = 7'h27 == io_i_rename_table_19 ? io_i_pregs_39 : _GEN_2470; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2472 = 7'h28 == io_i_rename_table_19 ? io_i_pregs_40 : _GEN_2471; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2473 = 7'h29 == io_i_rename_table_19 ? io_i_pregs_41 : _GEN_2472; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2474 = 7'h2a == io_i_rename_table_19 ? io_i_pregs_42 : _GEN_2473; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2475 = 7'h2b == io_i_rename_table_19 ? io_i_pregs_43 : _GEN_2474; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2476 = 7'h2c == io_i_rename_table_19 ? io_i_pregs_44 : _GEN_2475; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2477 = 7'h2d == io_i_rename_table_19 ? io_i_pregs_45 : _GEN_2476; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2478 = 7'h2e == io_i_rename_table_19 ? io_i_pregs_46 : _GEN_2477; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2479 = 7'h2f == io_i_rename_table_19 ? io_i_pregs_47 : _GEN_2478; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2480 = 7'h30 == io_i_rename_table_19 ? io_i_pregs_48 : _GEN_2479; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2481 = 7'h31 == io_i_rename_table_19 ? io_i_pregs_49 : _GEN_2480; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2482 = 7'h32 == io_i_rename_table_19 ? io_i_pregs_50 : _GEN_2481; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2483 = 7'h33 == io_i_rename_table_19 ? io_i_pregs_51 : _GEN_2482; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2484 = 7'h34 == io_i_rename_table_19 ? io_i_pregs_52 : _GEN_2483; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2485 = 7'h35 == io_i_rename_table_19 ? io_i_pregs_53 : _GEN_2484; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2486 = 7'h36 == io_i_rename_table_19 ? io_i_pregs_54 : _GEN_2485; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2487 = 7'h37 == io_i_rename_table_19 ? io_i_pregs_55 : _GEN_2486; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2488 = 7'h38 == io_i_rename_table_19 ? io_i_pregs_56 : _GEN_2487; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2489 = 7'h39 == io_i_rename_table_19 ? io_i_pregs_57 : _GEN_2488; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2490 = 7'h3a == io_i_rename_table_19 ? io_i_pregs_58 : _GEN_2489; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2491 = 7'h3b == io_i_rename_table_19 ? io_i_pregs_59 : _GEN_2490; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2492 = 7'h3c == io_i_rename_table_19 ? io_i_pregs_60 : _GEN_2491; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2493 = 7'h3d == io_i_rename_table_19 ? io_i_pregs_61 : _GEN_2492; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2494 = 7'h3e == io_i_rename_table_19 ? io_i_pregs_62 : _GEN_2493; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2495 = 7'h3f == io_i_rename_table_19 ? io_i_pregs_63 : _GEN_2494; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2496 = 7'h40 == io_i_rename_table_19 ? io_i_pregs_64 : _GEN_2495; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2497 = 7'h41 == io_i_rename_table_19 ? io_i_pregs_65 : _GEN_2496; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2498 = 7'h42 == io_i_rename_table_19 ? io_i_pregs_66 : _GEN_2497; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2499 = 7'h43 == io_i_rename_table_19 ? io_i_pregs_67 : _GEN_2498; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2500 = 7'h44 == io_i_rename_table_19 ? io_i_pregs_68 : _GEN_2499; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2501 = 7'h45 == io_i_rename_table_19 ? io_i_pregs_69 : _GEN_2500; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2502 = 7'h46 == io_i_rename_table_19 ? io_i_pregs_70 : _GEN_2501; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2503 = 7'h47 == io_i_rename_table_19 ? io_i_pregs_71 : _GEN_2502; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2504 = 7'h48 == io_i_rename_table_19 ? io_i_pregs_72 : _GEN_2503; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2505 = 7'h49 == io_i_rename_table_19 ? io_i_pregs_73 : _GEN_2504; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2506 = 7'h4a == io_i_rename_table_19 ? io_i_pregs_74 : _GEN_2505; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2507 = 7'h4b == io_i_rename_table_19 ? io_i_pregs_75 : _GEN_2506; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2508 = 7'h4c == io_i_rename_table_19 ? io_i_pregs_76 : _GEN_2507; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2509 = 7'h4d == io_i_rename_table_19 ? io_i_pregs_77 : _GEN_2508; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2510 = 7'h4e == io_i_rename_table_19 ? io_i_pregs_78 : _GEN_2509; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2511 = 7'h4f == io_i_rename_table_19 ? io_i_pregs_79 : _GEN_2510; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2512 = 7'h50 == io_i_rename_table_19 ? io_i_pregs_80 : _GEN_2511; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2513 = 7'h51 == io_i_rename_table_19 ? io_i_pregs_81 : _GEN_2512; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2514 = 7'h52 == io_i_rename_table_19 ? io_i_pregs_82 : _GEN_2513; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2515 = 7'h53 == io_i_rename_table_19 ? io_i_pregs_83 : _GEN_2514; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2516 = 7'h54 == io_i_rename_table_19 ? io_i_pregs_84 : _GEN_2515; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2517 = 7'h55 == io_i_rename_table_19 ? io_i_pregs_85 : _GEN_2516; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2518 = 7'h56 == io_i_rename_table_19 ? io_i_pregs_86 : _GEN_2517; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2519 = 7'h57 == io_i_rename_table_19 ? io_i_pregs_87 : _GEN_2518; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2520 = 7'h58 == io_i_rename_table_19 ? io_i_pregs_88 : _GEN_2519; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2521 = 7'h59 == io_i_rename_table_19 ? io_i_pregs_89 : _GEN_2520; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2522 = 7'h5a == io_i_rename_table_19 ? io_i_pregs_90 : _GEN_2521; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2523 = 7'h5b == io_i_rename_table_19 ? io_i_pregs_91 : _GEN_2522; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2524 = 7'h5c == io_i_rename_table_19 ? io_i_pregs_92 : _GEN_2523; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2525 = 7'h5d == io_i_rename_table_19 ? io_i_pregs_93 : _GEN_2524; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2526 = 7'h5e == io_i_rename_table_19 ? io_i_pregs_94 : _GEN_2525; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2527 = 7'h5f == io_i_rename_table_19 ? io_i_pregs_95 : _GEN_2526; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2528 = 7'h60 == io_i_rename_table_19 ? io_i_pregs_96 : _GEN_2527; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2529 = 7'h61 == io_i_rename_table_19 ? io_i_pregs_97 : _GEN_2528; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2530 = 7'h62 == io_i_rename_table_19 ? io_i_pregs_98 : _GEN_2529; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2531 = 7'h63 == io_i_rename_table_19 ? io_i_pregs_99 : _GEN_2530; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2532 = 7'h64 == io_i_rename_table_19 ? io_i_pregs_100 : _GEN_2531; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2533 = 7'h65 == io_i_rename_table_19 ? io_i_pregs_101 : _GEN_2532; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2534 = 7'h66 == io_i_rename_table_19 ? io_i_pregs_102 : _GEN_2533; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2535 = 7'h67 == io_i_rename_table_19 ? io_i_pregs_103 : _GEN_2534; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2536 = 7'h68 == io_i_rename_table_19 ? io_i_pregs_104 : _GEN_2535; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2537 = 7'h69 == io_i_rename_table_19 ? io_i_pregs_105 : _GEN_2536; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2538 = 7'h6a == io_i_rename_table_19 ? io_i_pregs_106 : _GEN_2537; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2539 = 7'h6b == io_i_rename_table_19 ? io_i_pregs_107 : _GEN_2538; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2540 = 7'h6c == io_i_rename_table_19 ? io_i_pregs_108 : _GEN_2539; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2541 = 7'h6d == io_i_rename_table_19 ? io_i_pregs_109 : _GEN_2540; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2542 = 7'h6e == io_i_rename_table_19 ? io_i_pregs_110 : _GEN_2541; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2543 = 7'h6f == io_i_rename_table_19 ? io_i_pregs_111 : _GEN_2542; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2544 = 7'h70 == io_i_rename_table_19 ? io_i_pregs_112 : _GEN_2543; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2545 = 7'h71 == io_i_rename_table_19 ? io_i_pregs_113 : _GEN_2544; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2546 = 7'h72 == io_i_rename_table_19 ? io_i_pregs_114 : _GEN_2545; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2547 = 7'h73 == io_i_rename_table_19 ? io_i_pregs_115 : _GEN_2546; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2548 = 7'h74 == io_i_rename_table_19 ? io_i_pregs_116 : _GEN_2547; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2549 = 7'h75 == io_i_rename_table_19 ? io_i_pregs_117 : _GEN_2548; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2550 = 7'h76 == io_i_rename_table_19 ? io_i_pregs_118 : _GEN_2549; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2551 = 7'h77 == io_i_rename_table_19 ? io_i_pregs_119 : _GEN_2550; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2552 = 7'h78 == io_i_rename_table_19 ? io_i_pregs_120 : _GEN_2551; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2553 = 7'h79 == io_i_rename_table_19 ? io_i_pregs_121 : _GEN_2552; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2554 = 7'h7a == io_i_rename_table_19 ? io_i_pregs_122 : _GEN_2553; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2555 = 7'h7b == io_i_rename_table_19 ? io_i_pregs_123 : _GEN_2554; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2556 = 7'h7c == io_i_rename_table_19 ? io_i_pregs_124 : _GEN_2555; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2557 = 7'h7d == io_i_rename_table_19 ? io_i_pregs_125 : _GEN_2556; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2558 = 7'h7e == io_i_rename_table_19 ? io_i_pregs_126 : _GEN_2557; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2561 = 7'h1 == io_i_rename_table_20 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2562 = 7'h2 == io_i_rename_table_20 ? io_i_pregs_2 : _GEN_2561; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2563 = 7'h3 == io_i_rename_table_20 ? io_i_pregs_3 : _GEN_2562; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2564 = 7'h4 == io_i_rename_table_20 ? io_i_pregs_4 : _GEN_2563; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2565 = 7'h5 == io_i_rename_table_20 ? io_i_pregs_5 : _GEN_2564; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2566 = 7'h6 == io_i_rename_table_20 ? io_i_pregs_6 : _GEN_2565; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2567 = 7'h7 == io_i_rename_table_20 ? io_i_pregs_7 : _GEN_2566; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2568 = 7'h8 == io_i_rename_table_20 ? io_i_pregs_8 : _GEN_2567; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2569 = 7'h9 == io_i_rename_table_20 ? io_i_pregs_9 : _GEN_2568; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2570 = 7'ha == io_i_rename_table_20 ? io_i_pregs_10 : _GEN_2569; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2571 = 7'hb == io_i_rename_table_20 ? io_i_pregs_11 : _GEN_2570; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2572 = 7'hc == io_i_rename_table_20 ? io_i_pregs_12 : _GEN_2571; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2573 = 7'hd == io_i_rename_table_20 ? io_i_pregs_13 : _GEN_2572; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2574 = 7'he == io_i_rename_table_20 ? io_i_pregs_14 : _GEN_2573; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2575 = 7'hf == io_i_rename_table_20 ? io_i_pregs_15 : _GEN_2574; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2576 = 7'h10 == io_i_rename_table_20 ? io_i_pregs_16 : _GEN_2575; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2577 = 7'h11 == io_i_rename_table_20 ? io_i_pregs_17 : _GEN_2576; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2578 = 7'h12 == io_i_rename_table_20 ? io_i_pregs_18 : _GEN_2577; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2579 = 7'h13 == io_i_rename_table_20 ? io_i_pregs_19 : _GEN_2578; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2580 = 7'h14 == io_i_rename_table_20 ? io_i_pregs_20 : _GEN_2579; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2581 = 7'h15 == io_i_rename_table_20 ? io_i_pregs_21 : _GEN_2580; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2582 = 7'h16 == io_i_rename_table_20 ? io_i_pregs_22 : _GEN_2581; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2583 = 7'h17 == io_i_rename_table_20 ? io_i_pregs_23 : _GEN_2582; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2584 = 7'h18 == io_i_rename_table_20 ? io_i_pregs_24 : _GEN_2583; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2585 = 7'h19 == io_i_rename_table_20 ? io_i_pregs_25 : _GEN_2584; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2586 = 7'h1a == io_i_rename_table_20 ? io_i_pregs_26 : _GEN_2585; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2587 = 7'h1b == io_i_rename_table_20 ? io_i_pregs_27 : _GEN_2586; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2588 = 7'h1c == io_i_rename_table_20 ? io_i_pregs_28 : _GEN_2587; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2589 = 7'h1d == io_i_rename_table_20 ? io_i_pregs_29 : _GEN_2588; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2590 = 7'h1e == io_i_rename_table_20 ? io_i_pregs_30 : _GEN_2589; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2591 = 7'h1f == io_i_rename_table_20 ? io_i_pregs_31 : _GEN_2590; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2592 = 7'h20 == io_i_rename_table_20 ? io_i_pregs_32 : _GEN_2591; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2593 = 7'h21 == io_i_rename_table_20 ? io_i_pregs_33 : _GEN_2592; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2594 = 7'h22 == io_i_rename_table_20 ? io_i_pregs_34 : _GEN_2593; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2595 = 7'h23 == io_i_rename_table_20 ? io_i_pregs_35 : _GEN_2594; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2596 = 7'h24 == io_i_rename_table_20 ? io_i_pregs_36 : _GEN_2595; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2597 = 7'h25 == io_i_rename_table_20 ? io_i_pregs_37 : _GEN_2596; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2598 = 7'h26 == io_i_rename_table_20 ? io_i_pregs_38 : _GEN_2597; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2599 = 7'h27 == io_i_rename_table_20 ? io_i_pregs_39 : _GEN_2598; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2600 = 7'h28 == io_i_rename_table_20 ? io_i_pregs_40 : _GEN_2599; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2601 = 7'h29 == io_i_rename_table_20 ? io_i_pregs_41 : _GEN_2600; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2602 = 7'h2a == io_i_rename_table_20 ? io_i_pregs_42 : _GEN_2601; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2603 = 7'h2b == io_i_rename_table_20 ? io_i_pregs_43 : _GEN_2602; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2604 = 7'h2c == io_i_rename_table_20 ? io_i_pregs_44 : _GEN_2603; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2605 = 7'h2d == io_i_rename_table_20 ? io_i_pregs_45 : _GEN_2604; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2606 = 7'h2e == io_i_rename_table_20 ? io_i_pregs_46 : _GEN_2605; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2607 = 7'h2f == io_i_rename_table_20 ? io_i_pregs_47 : _GEN_2606; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2608 = 7'h30 == io_i_rename_table_20 ? io_i_pregs_48 : _GEN_2607; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2609 = 7'h31 == io_i_rename_table_20 ? io_i_pregs_49 : _GEN_2608; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2610 = 7'h32 == io_i_rename_table_20 ? io_i_pregs_50 : _GEN_2609; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2611 = 7'h33 == io_i_rename_table_20 ? io_i_pregs_51 : _GEN_2610; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2612 = 7'h34 == io_i_rename_table_20 ? io_i_pregs_52 : _GEN_2611; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2613 = 7'h35 == io_i_rename_table_20 ? io_i_pregs_53 : _GEN_2612; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2614 = 7'h36 == io_i_rename_table_20 ? io_i_pregs_54 : _GEN_2613; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2615 = 7'h37 == io_i_rename_table_20 ? io_i_pregs_55 : _GEN_2614; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2616 = 7'h38 == io_i_rename_table_20 ? io_i_pregs_56 : _GEN_2615; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2617 = 7'h39 == io_i_rename_table_20 ? io_i_pregs_57 : _GEN_2616; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2618 = 7'h3a == io_i_rename_table_20 ? io_i_pregs_58 : _GEN_2617; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2619 = 7'h3b == io_i_rename_table_20 ? io_i_pregs_59 : _GEN_2618; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2620 = 7'h3c == io_i_rename_table_20 ? io_i_pregs_60 : _GEN_2619; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2621 = 7'h3d == io_i_rename_table_20 ? io_i_pregs_61 : _GEN_2620; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2622 = 7'h3e == io_i_rename_table_20 ? io_i_pregs_62 : _GEN_2621; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2623 = 7'h3f == io_i_rename_table_20 ? io_i_pregs_63 : _GEN_2622; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2624 = 7'h40 == io_i_rename_table_20 ? io_i_pregs_64 : _GEN_2623; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2625 = 7'h41 == io_i_rename_table_20 ? io_i_pregs_65 : _GEN_2624; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2626 = 7'h42 == io_i_rename_table_20 ? io_i_pregs_66 : _GEN_2625; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2627 = 7'h43 == io_i_rename_table_20 ? io_i_pregs_67 : _GEN_2626; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2628 = 7'h44 == io_i_rename_table_20 ? io_i_pregs_68 : _GEN_2627; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2629 = 7'h45 == io_i_rename_table_20 ? io_i_pregs_69 : _GEN_2628; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2630 = 7'h46 == io_i_rename_table_20 ? io_i_pregs_70 : _GEN_2629; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2631 = 7'h47 == io_i_rename_table_20 ? io_i_pregs_71 : _GEN_2630; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2632 = 7'h48 == io_i_rename_table_20 ? io_i_pregs_72 : _GEN_2631; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2633 = 7'h49 == io_i_rename_table_20 ? io_i_pregs_73 : _GEN_2632; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2634 = 7'h4a == io_i_rename_table_20 ? io_i_pregs_74 : _GEN_2633; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2635 = 7'h4b == io_i_rename_table_20 ? io_i_pregs_75 : _GEN_2634; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2636 = 7'h4c == io_i_rename_table_20 ? io_i_pregs_76 : _GEN_2635; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2637 = 7'h4d == io_i_rename_table_20 ? io_i_pregs_77 : _GEN_2636; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2638 = 7'h4e == io_i_rename_table_20 ? io_i_pregs_78 : _GEN_2637; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2639 = 7'h4f == io_i_rename_table_20 ? io_i_pregs_79 : _GEN_2638; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2640 = 7'h50 == io_i_rename_table_20 ? io_i_pregs_80 : _GEN_2639; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2641 = 7'h51 == io_i_rename_table_20 ? io_i_pregs_81 : _GEN_2640; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2642 = 7'h52 == io_i_rename_table_20 ? io_i_pregs_82 : _GEN_2641; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2643 = 7'h53 == io_i_rename_table_20 ? io_i_pregs_83 : _GEN_2642; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2644 = 7'h54 == io_i_rename_table_20 ? io_i_pregs_84 : _GEN_2643; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2645 = 7'h55 == io_i_rename_table_20 ? io_i_pregs_85 : _GEN_2644; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2646 = 7'h56 == io_i_rename_table_20 ? io_i_pregs_86 : _GEN_2645; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2647 = 7'h57 == io_i_rename_table_20 ? io_i_pregs_87 : _GEN_2646; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2648 = 7'h58 == io_i_rename_table_20 ? io_i_pregs_88 : _GEN_2647; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2649 = 7'h59 == io_i_rename_table_20 ? io_i_pregs_89 : _GEN_2648; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2650 = 7'h5a == io_i_rename_table_20 ? io_i_pregs_90 : _GEN_2649; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2651 = 7'h5b == io_i_rename_table_20 ? io_i_pregs_91 : _GEN_2650; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2652 = 7'h5c == io_i_rename_table_20 ? io_i_pregs_92 : _GEN_2651; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2653 = 7'h5d == io_i_rename_table_20 ? io_i_pregs_93 : _GEN_2652; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2654 = 7'h5e == io_i_rename_table_20 ? io_i_pregs_94 : _GEN_2653; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2655 = 7'h5f == io_i_rename_table_20 ? io_i_pregs_95 : _GEN_2654; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2656 = 7'h60 == io_i_rename_table_20 ? io_i_pregs_96 : _GEN_2655; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2657 = 7'h61 == io_i_rename_table_20 ? io_i_pregs_97 : _GEN_2656; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2658 = 7'h62 == io_i_rename_table_20 ? io_i_pregs_98 : _GEN_2657; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2659 = 7'h63 == io_i_rename_table_20 ? io_i_pregs_99 : _GEN_2658; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2660 = 7'h64 == io_i_rename_table_20 ? io_i_pregs_100 : _GEN_2659; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2661 = 7'h65 == io_i_rename_table_20 ? io_i_pregs_101 : _GEN_2660; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2662 = 7'h66 == io_i_rename_table_20 ? io_i_pregs_102 : _GEN_2661; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2663 = 7'h67 == io_i_rename_table_20 ? io_i_pregs_103 : _GEN_2662; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2664 = 7'h68 == io_i_rename_table_20 ? io_i_pregs_104 : _GEN_2663; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2665 = 7'h69 == io_i_rename_table_20 ? io_i_pregs_105 : _GEN_2664; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2666 = 7'h6a == io_i_rename_table_20 ? io_i_pregs_106 : _GEN_2665; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2667 = 7'h6b == io_i_rename_table_20 ? io_i_pregs_107 : _GEN_2666; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2668 = 7'h6c == io_i_rename_table_20 ? io_i_pregs_108 : _GEN_2667; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2669 = 7'h6d == io_i_rename_table_20 ? io_i_pregs_109 : _GEN_2668; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2670 = 7'h6e == io_i_rename_table_20 ? io_i_pregs_110 : _GEN_2669; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2671 = 7'h6f == io_i_rename_table_20 ? io_i_pregs_111 : _GEN_2670; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2672 = 7'h70 == io_i_rename_table_20 ? io_i_pregs_112 : _GEN_2671; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2673 = 7'h71 == io_i_rename_table_20 ? io_i_pregs_113 : _GEN_2672; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2674 = 7'h72 == io_i_rename_table_20 ? io_i_pregs_114 : _GEN_2673; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2675 = 7'h73 == io_i_rename_table_20 ? io_i_pregs_115 : _GEN_2674; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2676 = 7'h74 == io_i_rename_table_20 ? io_i_pregs_116 : _GEN_2675; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2677 = 7'h75 == io_i_rename_table_20 ? io_i_pregs_117 : _GEN_2676; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2678 = 7'h76 == io_i_rename_table_20 ? io_i_pregs_118 : _GEN_2677; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2679 = 7'h77 == io_i_rename_table_20 ? io_i_pregs_119 : _GEN_2678; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2680 = 7'h78 == io_i_rename_table_20 ? io_i_pregs_120 : _GEN_2679; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2681 = 7'h79 == io_i_rename_table_20 ? io_i_pregs_121 : _GEN_2680; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2682 = 7'h7a == io_i_rename_table_20 ? io_i_pregs_122 : _GEN_2681; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2683 = 7'h7b == io_i_rename_table_20 ? io_i_pregs_123 : _GEN_2682; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2684 = 7'h7c == io_i_rename_table_20 ? io_i_pregs_124 : _GEN_2683; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2685 = 7'h7d == io_i_rename_table_20 ? io_i_pregs_125 : _GEN_2684; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2686 = 7'h7e == io_i_rename_table_20 ? io_i_pregs_126 : _GEN_2685; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2689 = 7'h1 == io_i_rename_table_21 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2690 = 7'h2 == io_i_rename_table_21 ? io_i_pregs_2 : _GEN_2689; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2691 = 7'h3 == io_i_rename_table_21 ? io_i_pregs_3 : _GEN_2690; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2692 = 7'h4 == io_i_rename_table_21 ? io_i_pregs_4 : _GEN_2691; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2693 = 7'h5 == io_i_rename_table_21 ? io_i_pregs_5 : _GEN_2692; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2694 = 7'h6 == io_i_rename_table_21 ? io_i_pregs_6 : _GEN_2693; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2695 = 7'h7 == io_i_rename_table_21 ? io_i_pregs_7 : _GEN_2694; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2696 = 7'h8 == io_i_rename_table_21 ? io_i_pregs_8 : _GEN_2695; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2697 = 7'h9 == io_i_rename_table_21 ? io_i_pregs_9 : _GEN_2696; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2698 = 7'ha == io_i_rename_table_21 ? io_i_pregs_10 : _GEN_2697; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2699 = 7'hb == io_i_rename_table_21 ? io_i_pregs_11 : _GEN_2698; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2700 = 7'hc == io_i_rename_table_21 ? io_i_pregs_12 : _GEN_2699; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2701 = 7'hd == io_i_rename_table_21 ? io_i_pregs_13 : _GEN_2700; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2702 = 7'he == io_i_rename_table_21 ? io_i_pregs_14 : _GEN_2701; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2703 = 7'hf == io_i_rename_table_21 ? io_i_pregs_15 : _GEN_2702; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2704 = 7'h10 == io_i_rename_table_21 ? io_i_pregs_16 : _GEN_2703; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2705 = 7'h11 == io_i_rename_table_21 ? io_i_pregs_17 : _GEN_2704; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2706 = 7'h12 == io_i_rename_table_21 ? io_i_pregs_18 : _GEN_2705; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2707 = 7'h13 == io_i_rename_table_21 ? io_i_pregs_19 : _GEN_2706; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2708 = 7'h14 == io_i_rename_table_21 ? io_i_pregs_20 : _GEN_2707; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2709 = 7'h15 == io_i_rename_table_21 ? io_i_pregs_21 : _GEN_2708; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2710 = 7'h16 == io_i_rename_table_21 ? io_i_pregs_22 : _GEN_2709; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2711 = 7'h17 == io_i_rename_table_21 ? io_i_pregs_23 : _GEN_2710; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2712 = 7'h18 == io_i_rename_table_21 ? io_i_pregs_24 : _GEN_2711; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2713 = 7'h19 == io_i_rename_table_21 ? io_i_pregs_25 : _GEN_2712; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2714 = 7'h1a == io_i_rename_table_21 ? io_i_pregs_26 : _GEN_2713; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2715 = 7'h1b == io_i_rename_table_21 ? io_i_pregs_27 : _GEN_2714; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2716 = 7'h1c == io_i_rename_table_21 ? io_i_pregs_28 : _GEN_2715; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2717 = 7'h1d == io_i_rename_table_21 ? io_i_pregs_29 : _GEN_2716; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2718 = 7'h1e == io_i_rename_table_21 ? io_i_pregs_30 : _GEN_2717; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2719 = 7'h1f == io_i_rename_table_21 ? io_i_pregs_31 : _GEN_2718; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2720 = 7'h20 == io_i_rename_table_21 ? io_i_pregs_32 : _GEN_2719; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2721 = 7'h21 == io_i_rename_table_21 ? io_i_pregs_33 : _GEN_2720; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2722 = 7'h22 == io_i_rename_table_21 ? io_i_pregs_34 : _GEN_2721; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2723 = 7'h23 == io_i_rename_table_21 ? io_i_pregs_35 : _GEN_2722; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2724 = 7'h24 == io_i_rename_table_21 ? io_i_pregs_36 : _GEN_2723; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2725 = 7'h25 == io_i_rename_table_21 ? io_i_pregs_37 : _GEN_2724; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2726 = 7'h26 == io_i_rename_table_21 ? io_i_pregs_38 : _GEN_2725; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2727 = 7'h27 == io_i_rename_table_21 ? io_i_pregs_39 : _GEN_2726; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2728 = 7'h28 == io_i_rename_table_21 ? io_i_pregs_40 : _GEN_2727; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2729 = 7'h29 == io_i_rename_table_21 ? io_i_pregs_41 : _GEN_2728; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2730 = 7'h2a == io_i_rename_table_21 ? io_i_pregs_42 : _GEN_2729; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2731 = 7'h2b == io_i_rename_table_21 ? io_i_pregs_43 : _GEN_2730; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2732 = 7'h2c == io_i_rename_table_21 ? io_i_pregs_44 : _GEN_2731; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2733 = 7'h2d == io_i_rename_table_21 ? io_i_pregs_45 : _GEN_2732; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2734 = 7'h2e == io_i_rename_table_21 ? io_i_pregs_46 : _GEN_2733; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2735 = 7'h2f == io_i_rename_table_21 ? io_i_pregs_47 : _GEN_2734; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2736 = 7'h30 == io_i_rename_table_21 ? io_i_pregs_48 : _GEN_2735; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2737 = 7'h31 == io_i_rename_table_21 ? io_i_pregs_49 : _GEN_2736; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2738 = 7'h32 == io_i_rename_table_21 ? io_i_pregs_50 : _GEN_2737; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2739 = 7'h33 == io_i_rename_table_21 ? io_i_pregs_51 : _GEN_2738; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2740 = 7'h34 == io_i_rename_table_21 ? io_i_pregs_52 : _GEN_2739; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2741 = 7'h35 == io_i_rename_table_21 ? io_i_pregs_53 : _GEN_2740; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2742 = 7'h36 == io_i_rename_table_21 ? io_i_pregs_54 : _GEN_2741; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2743 = 7'h37 == io_i_rename_table_21 ? io_i_pregs_55 : _GEN_2742; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2744 = 7'h38 == io_i_rename_table_21 ? io_i_pregs_56 : _GEN_2743; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2745 = 7'h39 == io_i_rename_table_21 ? io_i_pregs_57 : _GEN_2744; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2746 = 7'h3a == io_i_rename_table_21 ? io_i_pregs_58 : _GEN_2745; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2747 = 7'h3b == io_i_rename_table_21 ? io_i_pregs_59 : _GEN_2746; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2748 = 7'h3c == io_i_rename_table_21 ? io_i_pregs_60 : _GEN_2747; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2749 = 7'h3d == io_i_rename_table_21 ? io_i_pregs_61 : _GEN_2748; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2750 = 7'h3e == io_i_rename_table_21 ? io_i_pregs_62 : _GEN_2749; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2751 = 7'h3f == io_i_rename_table_21 ? io_i_pregs_63 : _GEN_2750; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2752 = 7'h40 == io_i_rename_table_21 ? io_i_pregs_64 : _GEN_2751; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2753 = 7'h41 == io_i_rename_table_21 ? io_i_pregs_65 : _GEN_2752; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2754 = 7'h42 == io_i_rename_table_21 ? io_i_pregs_66 : _GEN_2753; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2755 = 7'h43 == io_i_rename_table_21 ? io_i_pregs_67 : _GEN_2754; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2756 = 7'h44 == io_i_rename_table_21 ? io_i_pregs_68 : _GEN_2755; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2757 = 7'h45 == io_i_rename_table_21 ? io_i_pregs_69 : _GEN_2756; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2758 = 7'h46 == io_i_rename_table_21 ? io_i_pregs_70 : _GEN_2757; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2759 = 7'h47 == io_i_rename_table_21 ? io_i_pregs_71 : _GEN_2758; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2760 = 7'h48 == io_i_rename_table_21 ? io_i_pregs_72 : _GEN_2759; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2761 = 7'h49 == io_i_rename_table_21 ? io_i_pregs_73 : _GEN_2760; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2762 = 7'h4a == io_i_rename_table_21 ? io_i_pregs_74 : _GEN_2761; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2763 = 7'h4b == io_i_rename_table_21 ? io_i_pregs_75 : _GEN_2762; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2764 = 7'h4c == io_i_rename_table_21 ? io_i_pregs_76 : _GEN_2763; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2765 = 7'h4d == io_i_rename_table_21 ? io_i_pregs_77 : _GEN_2764; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2766 = 7'h4e == io_i_rename_table_21 ? io_i_pregs_78 : _GEN_2765; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2767 = 7'h4f == io_i_rename_table_21 ? io_i_pregs_79 : _GEN_2766; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2768 = 7'h50 == io_i_rename_table_21 ? io_i_pregs_80 : _GEN_2767; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2769 = 7'h51 == io_i_rename_table_21 ? io_i_pregs_81 : _GEN_2768; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2770 = 7'h52 == io_i_rename_table_21 ? io_i_pregs_82 : _GEN_2769; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2771 = 7'h53 == io_i_rename_table_21 ? io_i_pregs_83 : _GEN_2770; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2772 = 7'h54 == io_i_rename_table_21 ? io_i_pregs_84 : _GEN_2771; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2773 = 7'h55 == io_i_rename_table_21 ? io_i_pregs_85 : _GEN_2772; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2774 = 7'h56 == io_i_rename_table_21 ? io_i_pregs_86 : _GEN_2773; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2775 = 7'h57 == io_i_rename_table_21 ? io_i_pregs_87 : _GEN_2774; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2776 = 7'h58 == io_i_rename_table_21 ? io_i_pregs_88 : _GEN_2775; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2777 = 7'h59 == io_i_rename_table_21 ? io_i_pregs_89 : _GEN_2776; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2778 = 7'h5a == io_i_rename_table_21 ? io_i_pregs_90 : _GEN_2777; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2779 = 7'h5b == io_i_rename_table_21 ? io_i_pregs_91 : _GEN_2778; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2780 = 7'h5c == io_i_rename_table_21 ? io_i_pregs_92 : _GEN_2779; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2781 = 7'h5d == io_i_rename_table_21 ? io_i_pregs_93 : _GEN_2780; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2782 = 7'h5e == io_i_rename_table_21 ? io_i_pregs_94 : _GEN_2781; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2783 = 7'h5f == io_i_rename_table_21 ? io_i_pregs_95 : _GEN_2782; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2784 = 7'h60 == io_i_rename_table_21 ? io_i_pregs_96 : _GEN_2783; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2785 = 7'h61 == io_i_rename_table_21 ? io_i_pregs_97 : _GEN_2784; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2786 = 7'h62 == io_i_rename_table_21 ? io_i_pregs_98 : _GEN_2785; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2787 = 7'h63 == io_i_rename_table_21 ? io_i_pregs_99 : _GEN_2786; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2788 = 7'h64 == io_i_rename_table_21 ? io_i_pregs_100 : _GEN_2787; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2789 = 7'h65 == io_i_rename_table_21 ? io_i_pregs_101 : _GEN_2788; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2790 = 7'h66 == io_i_rename_table_21 ? io_i_pregs_102 : _GEN_2789; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2791 = 7'h67 == io_i_rename_table_21 ? io_i_pregs_103 : _GEN_2790; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2792 = 7'h68 == io_i_rename_table_21 ? io_i_pregs_104 : _GEN_2791; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2793 = 7'h69 == io_i_rename_table_21 ? io_i_pregs_105 : _GEN_2792; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2794 = 7'h6a == io_i_rename_table_21 ? io_i_pregs_106 : _GEN_2793; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2795 = 7'h6b == io_i_rename_table_21 ? io_i_pregs_107 : _GEN_2794; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2796 = 7'h6c == io_i_rename_table_21 ? io_i_pregs_108 : _GEN_2795; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2797 = 7'h6d == io_i_rename_table_21 ? io_i_pregs_109 : _GEN_2796; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2798 = 7'h6e == io_i_rename_table_21 ? io_i_pregs_110 : _GEN_2797; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2799 = 7'h6f == io_i_rename_table_21 ? io_i_pregs_111 : _GEN_2798; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2800 = 7'h70 == io_i_rename_table_21 ? io_i_pregs_112 : _GEN_2799; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2801 = 7'h71 == io_i_rename_table_21 ? io_i_pregs_113 : _GEN_2800; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2802 = 7'h72 == io_i_rename_table_21 ? io_i_pregs_114 : _GEN_2801; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2803 = 7'h73 == io_i_rename_table_21 ? io_i_pregs_115 : _GEN_2802; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2804 = 7'h74 == io_i_rename_table_21 ? io_i_pregs_116 : _GEN_2803; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2805 = 7'h75 == io_i_rename_table_21 ? io_i_pregs_117 : _GEN_2804; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2806 = 7'h76 == io_i_rename_table_21 ? io_i_pregs_118 : _GEN_2805; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2807 = 7'h77 == io_i_rename_table_21 ? io_i_pregs_119 : _GEN_2806; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2808 = 7'h78 == io_i_rename_table_21 ? io_i_pregs_120 : _GEN_2807; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2809 = 7'h79 == io_i_rename_table_21 ? io_i_pregs_121 : _GEN_2808; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2810 = 7'h7a == io_i_rename_table_21 ? io_i_pregs_122 : _GEN_2809; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2811 = 7'h7b == io_i_rename_table_21 ? io_i_pregs_123 : _GEN_2810; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2812 = 7'h7c == io_i_rename_table_21 ? io_i_pregs_124 : _GEN_2811; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2813 = 7'h7d == io_i_rename_table_21 ? io_i_pregs_125 : _GEN_2812; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2814 = 7'h7e == io_i_rename_table_21 ? io_i_pregs_126 : _GEN_2813; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2817 = 7'h1 == io_i_rename_table_22 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2818 = 7'h2 == io_i_rename_table_22 ? io_i_pregs_2 : _GEN_2817; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2819 = 7'h3 == io_i_rename_table_22 ? io_i_pregs_3 : _GEN_2818; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2820 = 7'h4 == io_i_rename_table_22 ? io_i_pregs_4 : _GEN_2819; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2821 = 7'h5 == io_i_rename_table_22 ? io_i_pregs_5 : _GEN_2820; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2822 = 7'h6 == io_i_rename_table_22 ? io_i_pregs_6 : _GEN_2821; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2823 = 7'h7 == io_i_rename_table_22 ? io_i_pregs_7 : _GEN_2822; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2824 = 7'h8 == io_i_rename_table_22 ? io_i_pregs_8 : _GEN_2823; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2825 = 7'h9 == io_i_rename_table_22 ? io_i_pregs_9 : _GEN_2824; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2826 = 7'ha == io_i_rename_table_22 ? io_i_pregs_10 : _GEN_2825; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2827 = 7'hb == io_i_rename_table_22 ? io_i_pregs_11 : _GEN_2826; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2828 = 7'hc == io_i_rename_table_22 ? io_i_pregs_12 : _GEN_2827; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2829 = 7'hd == io_i_rename_table_22 ? io_i_pregs_13 : _GEN_2828; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2830 = 7'he == io_i_rename_table_22 ? io_i_pregs_14 : _GEN_2829; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2831 = 7'hf == io_i_rename_table_22 ? io_i_pregs_15 : _GEN_2830; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2832 = 7'h10 == io_i_rename_table_22 ? io_i_pregs_16 : _GEN_2831; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2833 = 7'h11 == io_i_rename_table_22 ? io_i_pregs_17 : _GEN_2832; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2834 = 7'h12 == io_i_rename_table_22 ? io_i_pregs_18 : _GEN_2833; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2835 = 7'h13 == io_i_rename_table_22 ? io_i_pregs_19 : _GEN_2834; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2836 = 7'h14 == io_i_rename_table_22 ? io_i_pregs_20 : _GEN_2835; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2837 = 7'h15 == io_i_rename_table_22 ? io_i_pregs_21 : _GEN_2836; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2838 = 7'h16 == io_i_rename_table_22 ? io_i_pregs_22 : _GEN_2837; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2839 = 7'h17 == io_i_rename_table_22 ? io_i_pregs_23 : _GEN_2838; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2840 = 7'h18 == io_i_rename_table_22 ? io_i_pregs_24 : _GEN_2839; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2841 = 7'h19 == io_i_rename_table_22 ? io_i_pregs_25 : _GEN_2840; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2842 = 7'h1a == io_i_rename_table_22 ? io_i_pregs_26 : _GEN_2841; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2843 = 7'h1b == io_i_rename_table_22 ? io_i_pregs_27 : _GEN_2842; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2844 = 7'h1c == io_i_rename_table_22 ? io_i_pregs_28 : _GEN_2843; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2845 = 7'h1d == io_i_rename_table_22 ? io_i_pregs_29 : _GEN_2844; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2846 = 7'h1e == io_i_rename_table_22 ? io_i_pregs_30 : _GEN_2845; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2847 = 7'h1f == io_i_rename_table_22 ? io_i_pregs_31 : _GEN_2846; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2848 = 7'h20 == io_i_rename_table_22 ? io_i_pregs_32 : _GEN_2847; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2849 = 7'h21 == io_i_rename_table_22 ? io_i_pregs_33 : _GEN_2848; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2850 = 7'h22 == io_i_rename_table_22 ? io_i_pregs_34 : _GEN_2849; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2851 = 7'h23 == io_i_rename_table_22 ? io_i_pregs_35 : _GEN_2850; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2852 = 7'h24 == io_i_rename_table_22 ? io_i_pregs_36 : _GEN_2851; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2853 = 7'h25 == io_i_rename_table_22 ? io_i_pregs_37 : _GEN_2852; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2854 = 7'h26 == io_i_rename_table_22 ? io_i_pregs_38 : _GEN_2853; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2855 = 7'h27 == io_i_rename_table_22 ? io_i_pregs_39 : _GEN_2854; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2856 = 7'h28 == io_i_rename_table_22 ? io_i_pregs_40 : _GEN_2855; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2857 = 7'h29 == io_i_rename_table_22 ? io_i_pregs_41 : _GEN_2856; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2858 = 7'h2a == io_i_rename_table_22 ? io_i_pregs_42 : _GEN_2857; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2859 = 7'h2b == io_i_rename_table_22 ? io_i_pregs_43 : _GEN_2858; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2860 = 7'h2c == io_i_rename_table_22 ? io_i_pregs_44 : _GEN_2859; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2861 = 7'h2d == io_i_rename_table_22 ? io_i_pregs_45 : _GEN_2860; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2862 = 7'h2e == io_i_rename_table_22 ? io_i_pregs_46 : _GEN_2861; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2863 = 7'h2f == io_i_rename_table_22 ? io_i_pregs_47 : _GEN_2862; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2864 = 7'h30 == io_i_rename_table_22 ? io_i_pregs_48 : _GEN_2863; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2865 = 7'h31 == io_i_rename_table_22 ? io_i_pregs_49 : _GEN_2864; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2866 = 7'h32 == io_i_rename_table_22 ? io_i_pregs_50 : _GEN_2865; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2867 = 7'h33 == io_i_rename_table_22 ? io_i_pregs_51 : _GEN_2866; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2868 = 7'h34 == io_i_rename_table_22 ? io_i_pregs_52 : _GEN_2867; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2869 = 7'h35 == io_i_rename_table_22 ? io_i_pregs_53 : _GEN_2868; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2870 = 7'h36 == io_i_rename_table_22 ? io_i_pregs_54 : _GEN_2869; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2871 = 7'h37 == io_i_rename_table_22 ? io_i_pregs_55 : _GEN_2870; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2872 = 7'h38 == io_i_rename_table_22 ? io_i_pregs_56 : _GEN_2871; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2873 = 7'h39 == io_i_rename_table_22 ? io_i_pregs_57 : _GEN_2872; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2874 = 7'h3a == io_i_rename_table_22 ? io_i_pregs_58 : _GEN_2873; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2875 = 7'h3b == io_i_rename_table_22 ? io_i_pregs_59 : _GEN_2874; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2876 = 7'h3c == io_i_rename_table_22 ? io_i_pregs_60 : _GEN_2875; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2877 = 7'h3d == io_i_rename_table_22 ? io_i_pregs_61 : _GEN_2876; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2878 = 7'h3e == io_i_rename_table_22 ? io_i_pregs_62 : _GEN_2877; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2879 = 7'h3f == io_i_rename_table_22 ? io_i_pregs_63 : _GEN_2878; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2880 = 7'h40 == io_i_rename_table_22 ? io_i_pregs_64 : _GEN_2879; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2881 = 7'h41 == io_i_rename_table_22 ? io_i_pregs_65 : _GEN_2880; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2882 = 7'h42 == io_i_rename_table_22 ? io_i_pregs_66 : _GEN_2881; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2883 = 7'h43 == io_i_rename_table_22 ? io_i_pregs_67 : _GEN_2882; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2884 = 7'h44 == io_i_rename_table_22 ? io_i_pregs_68 : _GEN_2883; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2885 = 7'h45 == io_i_rename_table_22 ? io_i_pregs_69 : _GEN_2884; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2886 = 7'h46 == io_i_rename_table_22 ? io_i_pregs_70 : _GEN_2885; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2887 = 7'h47 == io_i_rename_table_22 ? io_i_pregs_71 : _GEN_2886; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2888 = 7'h48 == io_i_rename_table_22 ? io_i_pregs_72 : _GEN_2887; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2889 = 7'h49 == io_i_rename_table_22 ? io_i_pregs_73 : _GEN_2888; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2890 = 7'h4a == io_i_rename_table_22 ? io_i_pregs_74 : _GEN_2889; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2891 = 7'h4b == io_i_rename_table_22 ? io_i_pregs_75 : _GEN_2890; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2892 = 7'h4c == io_i_rename_table_22 ? io_i_pregs_76 : _GEN_2891; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2893 = 7'h4d == io_i_rename_table_22 ? io_i_pregs_77 : _GEN_2892; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2894 = 7'h4e == io_i_rename_table_22 ? io_i_pregs_78 : _GEN_2893; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2895 = 7'h4f == io_i_rename_table_22 ? io_i_pregs_79 : _GEN_2894; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2896 = 7'h50 == io_i_rename_table_22 ? io_i_pregs_80 : _GEN_2895; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2897 = 7'h51 == io_i_rename_table_22 ? io_i_pregs_81 : _GEN_2896; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2898 = 7'h52 == io_i_rename_table_22 ? io_i_pregs_82 : _GEN_2897; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2899 = 7'h53 == io_i_rename_table_22 ? io_i_pregs_83 : _GEN_2898; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2900 = 7'h54 == io_i_rename_table_22 ? io_i_pregs_84 : _GEN_2899; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2901 = 7'h55 == io_i_rename_table_22 ? io_i_pregs_85 : _GEN_2900; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2902 = 7'h56 == io_i_rename_table_22 ? io_i_pregs_86 : _GEN_2901; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2903 = 7'h57 == io_i_rename_table_22 ? io_i_pregs_87 : _GEN_2902; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2904 = 7'h58 == io_i_rename_table_22 ? io_i_pregs_88 : _GEN_2903; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2905 = 7'h59 == io_i_rename_table_22 ? io_i_pregs_89 : _GEN_2904; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2906 = 7'h5a == io_i_rename_table_22 ? io_i_pregs_90 : _GEN_2905; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2907 = 7'h5b == io_i_rename_table_22 ? io_i_pregs_91 : _GEN_2906; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2908 = 7'h5c == io_i_rename_table_22 ? io_i_pregs_92 : _GEN_2907; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2909 = 7'h5d == io_i_rename_table_22 ? io_i_pregs_93 : _GEN_2908; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2910 = 7'h5e == io_i_rename_table_22 ? io_i_pregs_94 : _GEN_2909; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2911 = 7'h5f == io_i_rename_table_22 ? io_i_pregs_95 : _GEN_2910; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2912 = 7'h60 == io_i_rename_table_22 ? io_i_pregs_96 : _GEN_2911; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2913 = 7'h61 == io_i_rename_table_22 ? io_i_pregs_97 : _GEN_2912; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2914 = 7'h62 == io_i_rename_table_22 ? io_i_pregs_98 : _GEN_2913; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2915 = 7'h63 == io_i_rename_table_22 ? io_i_pregs_99 : _GEN_2914; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2916 = 7'h64 == io_i_rename_table_22 ? io_i_pregs_100 : _GEN_2915; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2917 = 7'h65 == io_i_rename_table_22 ? io_i_pregs_101 : _GEN_2916; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2918 = 7'h66 == io_i_rename_table_22 ? io_i_pregs_102 : _GEN_2917; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2919 = 7'h67 == io_i_rename_table_22 ? io_i_pregs_103 : _GEN_2918; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2920 = 7'h68 == io_i_rename_table_22 ? io_i_pregs_104 : _GEN_2919; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2921 = 7'h69 == io_i_rename_table_22 ? io_i_pregs_105 : _GEN_2920; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2922 = 7'h6a == io_i_rename_table_22 ? io_i_pregs_106 : _GEN_2921; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2923 = 7'h6b == io_i_rename_table_22 ? io_i_pregs_107 : _GEN_2922; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2924 = 7'h6c == io_i_rename_table_22 ? io_i_pregs_108 : _GEN_2923; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2925 = 7'h6d == io_i_rename_table_22 ? io_i_pregs_109 : _GEN_2924; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2926 = 7'h6e == io_i_rename_table_22 ? io_i_pregs_110 : _GEN_2925; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2927 = 7'h6f == io_i_rename_table_22 ? io_i_pregs_111 : _GEN_2926; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2928 = 7'h70 == io_i_rename_table_22 ? io_i_pregs_112 : _GEN_2927; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2929 = 7'h71 == io_i_rename_table_22 ? io_i_pregs_113 : _GEN_2928; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2930 = 7'h72 == io_i_rename_table_22 ? io_i_pregs_114 : _GEN_2929; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2931 = 7'h73 == io_i_rename_table_22 ? io_i_pregs_115 : _GEN_2930; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2932 = 7'h74 == io_i_rename_table_22 ? io_i_pregs_116 : _GEN_2931; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2933 = 7'h75 == io_i_rename_table_22 ? io_i_pregs_117 : _GEN_2932; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2934 = 7'h76 == io_i_rename_table_22 ? io_i_pregs_118 : _GEN_2933; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2935 = 7'h77 == io_i_rename_table_22 ? io_i_pregs_119 : _GEN_2934; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2936 = 7'h78 == io_i_rename_table_22 ? io_i_pregs_120 : _GEN_2935; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2937 = 7'h79 == io_i_rename_table_22 ? io_i_pregs_121 : _GEN_2936; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2938 = 7'h7a == io_i_rename_table_22 ? io_i_pregs_122 : _GEN_2937; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2939 = 7'h7b == io_i_rename_table_22 ? io_i_pregs_123 : _GEN_2938; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2940 = 7'h7c == io_i_rename_table_22 ? io_i_pregs_124 : _GEN_2939; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2941 = 7'h7d == io_i_rename_table_22 ? io_i_pregs_125 : _GEN_2940; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2942 = 7'h7e == io_i_rename_table_22 ? io_i_pregs_126 : _GEN_2941; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2945 = 7'h1 == io_i_rename_table_23 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2946 = 7'h2 == io_i_rename_table_23 ? io_i_pregs_2 : _GEN_2945; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2947 = 7'h3 == io_i_rename_table_23 ? io_i_pregs_3 : _GEN_2946; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2948 = 7'h4 == io_i_rename_table_23 ? io_i_pregs_4 : _GEN_2947; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2949 = 7'h5 == io_i_rename_table_23 ? io_i_pregs_5 : _GEN_2948; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2950 = 7'h6 == io_i_rename_table_23 ? io_i_pregs_6 : _GEN_2949; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2951 = 7'h7 == io_i_rename_table_23 ? io_i_pregs_7 : _GEN_2950; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2952 = 7'h8 == io_i_rename_table_23 ? io_i_pregs_8 : _GEN_2951; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2953 = 7'h9 == io_i_rename_table_23 ? io_i_pregs_9 : _GEN_2952; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2954 = 7'ha == io_i_rename_table_23 ? io_i_pregs_10 : _GEN_2953; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2955 = 7'hb == io_i_rename_table_23 ? io_i_pregs_11 : _GEN_2954; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2956 = 7'hc == io_i_rename_table_23 ? io_i_pregs_12 : _GEN_2955; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2957 = 7'hd == io_i_rename_table_23 ? io_i_pregs_13 : _GEN_2956; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2958 = 7'he == io_i_rename_table_23 ? io_i_pregs_14 : _GEN_2957; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2959 = 7'hf == io_i_rename_table_23 ? io_i_pregs_15 : _GEN_2958; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2960 = 7'h10 == io_i_rename_table_23 ? io_i_pregs_16 : _GEN_2959; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2961 = 7'h11 == io_i_rename_table_23 ? io_i_pregs_17 : _GEN_2960; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2962 = 7'h12 == io_i_rename_table_23 ? io_i_pregs_18 : _GEN_2961; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2963 = 7'h13 == io_i_rename_table_23 ? io_i_pregs_19 : _GEN_2962; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2964 = 7'h14 == io_i_rename_table_23 ? io_i_pregs_20 : _GEN_2963; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2965 = 7'h15 == io_i_rename_table_23 ? io_i_pregs_21 : _GEN_2964; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2966 = 7'h16 == io_i_rename_table_23 ? io_i_pregs_22 : _GEN_2965; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2967 = 7'h17 == io_i_rename_table_23 ? io_i_pregs_23 : _GEN_2966; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2968 = 7'h18 == io_i_rename_table_23 ? io_i_pregs_24 : _GEN_2967; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2969 = 7'h19 == io_i_rename_table_23 ? io_i_pregs_25 : _GEN_2968; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2970 = 7'h1a == io_i_rename_table_23 ? io_i_pregs_26 : _GEN_2969; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2971 = 7'h1b == io_i_rename_table_23 ? io_i_pregs_27 : _GEN_2970; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2972 = 7'h1c == io_i_rename_table_23 ? io_i_pregs_28 : _GEN_2971; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2973 = 7'h1d == io_i_rename_table_23 ? io_i_pregs_29 : _GEN_2972; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2974 = 7'h1e == io_i_rename_table_23 ? io_i_pregs_30 : _GEN_2973; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2975 = 7'h1f == io_i_rename_table_23 ? io_i_pregs_31 : _GEN_2974; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2976 = 7'h20 == io_i_rename_table_23 ? io_i_pregs_32 : _GEN_2975; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2977 = 7'h21 == io_i_rename_table_23 ? io_i_pregs_33 : _GEN_2976; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2978 = 7'h22 == io_i_rename_table_23 ? io_i_pregs_34 : _GEN_2977; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2979 = 7'h23 == io_i_rename_table_23 ? io_i_pregs_35 : _GEN_2978; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2980 = 7'h24 == io_i_rename_table_23 ? io_i_pregs_36 : _GEN_2979; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2981 = 7'h25 == io_i_rename_table_23 ? io_i_pregs_37 : _GEN_2980; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2982 = 7'h26 == io_i_rename_table_23 ? io_i_pregs_38 : _GEN_2981; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2983 = 7'h27 == io_i_rename_table_23 ? io_i_pregs_39 : _GEN_2982; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2984 = 7'h28 == io_i_rename_table_23 ? io_i_pregs_40 : _GEN_2983; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2985 = 7'h29 == io_i_rename_table_23 ? io_i_pregs_41 : _GEN_2984; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2986 = 7'h2a == io_i_rename_table_23 ? io_i_pregs_42 : _GEN_2985; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2987 = 7'h2b == io_i_rename_table_23 ? io_i_pregs_43 : _GEN_2986; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2988 = 7'h2c == io_i_rename_table_23 ? io_i_pregs_44 : _GEN_2987; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2989 = 7'h2d == io_i_rename_table_23 ? io_i_pregs_45 : _GEN_2988; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2990 = 7'h2e == io_i_rename_table_23 ? io_i_pregs_46 : _GEN_2989; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2991 = 7'h2f == io_i_rename_table_23 ? io_i_pregs_47 : _GEN_2990; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2992 = 7'h30 == io_i_rename_table_23 ? io_i_pregs_48 : _GEN_2991; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2993 = 7'h31 == io_i_rename_table_23 ? io_i_pregs_49 : _GEN_2992; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2994 = 7'h32 == io_i_rename_table_23 ? io_i_pregs_50 : _GEN_2993; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2995 = 7'h33 == io_i_rename_table_23 ? io_i_pregs_51 : _GEN_2994; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2996 = 7'h34 == io_i_rename_table_23 ? io_i_pregs_52 : _GEN_2995; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2997 = 7'h35 == io_i_rename_table_23 ? io_i_pregs_53 : _GEN_2996; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2998 = 7'h36 == io_i_rename_table_23 ? io_i_pregs_54 : _GEN_2997; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_2999 = 7'h37 == io_i_rename_table_23 ? io_i_pregs_55 : _GEN_2998; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3000 = 7'h38 == io_i_rename_table_23 ? io_i_pregs_56 : _GEN_2999; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3001 = 7'h39 == io_i_rename_table_23 ? io_i_pregs_57 : _GEN_3000; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3002 = 7'h3a == io_i_rename_table_23 ? io_i_pregs_58 : _GEN_3001; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3003 = 7'h3b == io_i_rename_table_23 ? io_i_pregs_59 : _GEN_3002; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3004 = 7'h3c == io_i_rename_table_23 ? io_i_pregs_60 : _GEN_3003; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3005 = 7'h3d == io_i_rename_table_23 ? io_i_pregs_61 : _GEN_3004; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3006 = 7'h3e == io_i_rename_table_23 ? io_i_pregs_62 : _GEN_3005; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3007 = 7'h3f == io_i_rename_table_23 ? io_i_pregs_63 : _GEN_3006; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3008 = 7'h40 == io_i_rename_table_23 ? io_i_pregs_64 : _GEN_3007; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3009 = 7'h41 == io_i_rename_table_23 ? io_i_pregs_65 : _GEN_3008; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3010 = 7'h42 == io_i_rename_table_23 ? io_i_pregs_66 : _GEN_3009; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3011 = 7'h43 == io_i_rename_table_23 ? io_i_pregs_67 : _GEN_3010; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3012 = 7'h44 == io_i_rename_table_23 ? io_i_pregs_68 : _GEN_3011; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3013 = 7'h45 == io_i_rename_table_23 ? io_i_pregs_69 : _GEN_3012; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3014 = 7'h46 == io_i_rename_table_23 ? io_i_pregs_70 : _GEN_3013; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3015 = 7'h47 == io_i_rename_table_23 ? io_i_pregs_71 : _GEN_3014; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3016 = 7'h48 == io_i_rename_table_23 ? io_i_pregs_72 : _GEN_3015; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3017 = 7'h49 == io_i_rename_table_23 ? io_i_pregs_73 : _GEN_3016; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3018 = 7'h4a == io_i_rename_table_23 ? io_i_pregs_74 : _GEN_3017; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3019 = 7'h4b == io_i_rename_table_23 ? io_i_pregs_75 : _GEN_3018; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3020 = 7'h4c == io_i_rename_table_23 ? io_i_pregs_76 : _GEN_3019; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3021 = 7'h4d == io_i_rename_table_23 ? io_i_pregs_77 : _GEN_3020; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3022 = 7'h4e == io_i_rename_table_23 ? io_i_pregs_78 : _GEN_3021; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3023 = 7'h4f == io_i_rename_table_23 ? io_i_pregs_79 : _GEN_3022; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3024 = 7'h50 == io_i_rename_table_23 ? io_i_pregs_80 : _GEN_3023; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3025 = 7'h51 == io_i_rename_table_23 ? io_i_pregs_81 : _GEN_3024; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3026 = 7'h52 == io_i_rename_table_23 ? io_i_pregs_82 : _GEN_3025; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3027 = 7'h53 == io_i_rename_table_23 ? io_i_pregs_83 : _GEN_3026; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3028 = 7'h54 == io_i_rename_table_23 ? io_i_pregs_84 : _GEN_3027; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3029 = 7'h55 == io_i_rename_table_23 ? io_i_pregs_85 : _GEN_3028; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3030 = 7'h56 == io_i_rename_table_23 ? io_i_pregs_86 : _GEN_3029; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3031 = 7'h57 == io_i_rename_table_23 ? io_i_pregs_87 : _GEN_3030; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3032 = 7'h58 == io_i_rename_table_23 ? io_i_pregs_88 : _GEN_3031; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3033 = 7'h59 == io_i_rename_table_23 ? io_i_pregs_89 : _GEN_3032; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3034 = 7'h5a == io_i_rename_table_23 ? io_i_pregs_90 : _GEN_3033; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3035 = 7'h5b == io_i_rename_table_23 ? io_i_pregs_91 : _GEN_3034; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3036 = 7'h5c == io_i_rename_table_23 ? io_i_pregs_92 : _GEN_3035; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3037 = 7'h5d == io_i_rename_table_23 ? io_i_pregs_93 : _GEN_3036; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3038 = 7'h5e == io_i_rename_table_23 ? io_i_pregs_94 : _GEN_3037; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3039 = 7'h5f == io_i_rename_table_23 ? io_i_pregs_95 : _GEN_3038; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3040 = 7'h60 == io_i_rename_table_23 ? io_i_pregs_96 : _GEN_3039; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3041 = 7'h61 == io_i_rename_table_23 ? io_i_pregs_97 : _GEN_3040; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3042 = 7'h62 == io_i_rename_table_23 ? io_i_pregs_98 : _GEN_3041; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3043 = 7'h63 == io_i_rename_table_23 ? io_i_pregs_99 : _GEN_3042; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3044 = 7'h64 == io_i_rename_table_23 ? io_i_pregs_100 : _GEN_3043; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3045 = 7'h65 == io_i_rename_table_23 ? io_i_pregs_101 : _GEN_3044; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3046 = 7'h66 == io_i_rename_table_23 ? io_i_pregs_102 : _GEN_3045; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3047 = 7'h67 == io_i_rename_table_23 ? io_i_pregs_103 : _GEN_3046; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3048 = 7'h68 == io_i_rename_table_23 ? io_i_pregs_104 : _GEN_3047; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3049 = 7'h69 == io_i_rename_table_23 ? io_i_pregs_105 : _GEN_3048; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3050 = 7'h6a == io_i_rename_table_23 ? io_i_pregs_106 : _GEN_3049; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3051 = 7'h6b == io_i_rename_table_23 ? io_i_pregs_107 : _GEN_3050; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3052 = 7'h6c == io_i_rename_table_23 ? io_i_pregs_108 : _GEN_3051; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3053 = 7'h6d == io_i_rename_table_23 ? io_i_pregs_109 : _GEN_3052; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3054 = 7'h6e == io_i_rename_table_23 ? io_i_pregs_110 : _GEN_3053; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3055 = 7'h6f == io_i_rename_table_23 ? io_i_pregs_111 : _GEN_3054; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3056 = 7'h70 == io_i_rename_table_23 ? io_i_pregs_112 : _GEN_3055; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3057 = 7'h71 == io_i_rename_table_23 ? io_i_pregs_113 : _GEN_3056; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3058 = 7'h72 == io_i_rename_table_23 ? io_i_pregs_114 : _GEN_3057; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3059 = 7'h73 == io_i_rename_table_23 ? io_i_pregs_115 : _GEN_3058; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3060 = 7'h74 == io_i_rename_table_23 ? io_i_pregs_116 : _GEN_3059; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3061 = 7'h75 == io_i_rename_table_23 ? io_i_pregs_117 : _GEN_3060; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3062 = 7'h76 == io_i_rename_table_23 ? io_i_pregs_118 : _GEN_3061; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3063 = 7'h77 == io_i_rename_table_23 ? io_i_pregs_119 : _GEN_3062; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3064 = 7'h78 == io_i_rename_table_23 ? io_i_pregs_120 : _GEN_3063; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3065 = 7'h79 == io_i_rename_table_23 ? io_i_pregs_121 : _GEN_3064; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3066 = 7'h7a == io_i_rename_table_23 ? io_i_pregs_122 : _GEN_3065; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3067 = 7'h7b == io_i_rename_table_23 ? io_i_pregs_123 : _GEN_3066; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3068 = 7'h7c == io_i_rename_table_23 ? io_i_pregs_124 : _GEN_3067; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3069 = 7'h7d == io_i_rename_table_23 ? io_i_pregs_125 : _GEN_3068; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3070 = 7'h7e == io_i_rename_table_23 ? io_i_pregs_126 : _GEN_3069; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3073 = 7'h1 == io_i_rename_table_24 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3074 = 7'h2 == io_i_rename_table_24 ? io_i_pregs_2 : _GEN_3073; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3075 = 7'h3 == io_i_rename_table_24 ? io_i_pregs_3 : _GEN_3074; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3076 = 7'h4 == io_i_rename_table_24 ? io_i_pregs_4 : _GEN_3075; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3077 = 7'h5 == io_i_rename_table_24 ? io_i_pregs_5 : _GEN_3076; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3078 = 7'h6 == io_i_rename_table_24 ? io_i_pregs_6 : _GEN_3077; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3079 = 7'h7 == io_i_rename_table_24 ? io_i_pregs_7 : _GEN_3078; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3080 = 7'h8 == io_i_rename_table_24 ? io_i_pregs_8 : _GEN_3079; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3081 = 7'h9 == io_i_rename_table_24 ? io_i_pregs_9 : _GEN_3080; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3082 = 7'ha == io_i_rename_table_24 ? io_i_pregs_10 : _GEN_3081; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3083 = 7'hb == io_i_rename_table_24 ? io_i_pregs_11 : _GEN_3082; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3084 = 7'hc == io_i_rename_table_24 ? io_i_pregs_12 : _GEN_3083; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3085 = 7'hd == io_i_rename_table_24 ? io_i_pregs_13 : _GEN_3084; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3086 = 7'he == io_i_rename_table_24 ? io_i_pregs_14 : _GEN_3085; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3087 = 7'hf == io_i_rename_table_24 ? io_i_pregs_15 : _GEN_3086; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3088 = 7'h10 == io_i_rename_table_24 ? io_i_pregs_16 : _GEN_3087; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3089 = 7'h11 == io_i_rename_table_24 ? io_i_pregs_17 : _GEN_3088; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3090 = 7'h12 == io_i_rename_table_24 ? io_i_pregs_18 : _GEN_3089; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3091 = 7'h13 == io_i_rename_table_24 ? io_i_pregs_19 : _GEN_3090; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3092 = 7'h14 == io_i_rename_table_24 ? io_i_pregs_20 : _GEN_3091; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3093 = 7'h15 == io_i_rename_table_24 ? io_i_pregs_21 : _GEN_3092; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3094 = 7'h16 == io_i_rename_table_24 ? io_i_pregs_22 : _GEN_3093; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3095 = 7'h17 == io_i_rename_table_24 ? io_i_pregs_23 : _GEN_3094; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3096 = 7'h18 == io_i_rename_table_24 ? io_i_pregs_24 : _GEN_3095; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3097 = 7'h19 == io_i_rename_table_24 ? io_i_pregs_25 : _GEN_3096; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3098 = 7'h1a == io_i_rename_table_24 ? io_i_pregs_26 : _GEN_3097; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3099 = 7'h1b == io_i_rename_table_24 ? io_i_pregs_27 : _GEN_3098; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3100 = 7'h1c == io_i_rename_table_24 ? io_i_pregs_28 : _GEN_3099; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3101 = 7'h1d == io_i_rename_table_24 ? io_i_pregs_29 : _GEN_3100; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3102 = 7'h1e == io_i_rename_table_24 ? io_i_pregs_30 : _GEN_3101; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3103 = 7'h1f == io_i_rename_table_24 ? io_i_pregs_31 : _GEN_3102; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3104 = 7'h20 == io_i_rename_table_24 ? io_i_pregs_32 : _GEN_3103; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3105 = 7'h21 == io_i_rename_table_24 ? io_i_pregs_33 : _GEN_3104; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3106 = 7'h22 == io_i_rename_table_24 ? io_i_pregs_34 : _GEN_3105; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3107 = 7'h23 == io_i_rename_table_24 ? io_i_pregs_35 : _GEN_3106; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3108 = 7'h24 == io_i_rename_table_24 ? io_i_pregs_36 : _GEN_3107; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3109 = 7'h25 == io_i_rename_table_24 ? io_i_pregs_37 : _GEN_3108; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3110 = 7'h26 == io_i_rename_table_24 ? io_i_pregs_38 : _GEN_3109; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3111 = 7'h27 == io_i_rename_table_24 ? io_i_pregs_39 : _GEN_3110; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3112 = 7'h28 == io_i_rename_table_24 ? io_i_pregs_40 : _GEN_3111; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3113 = 7'h29 == io_i_rename_table_24 ? io_i_pregs_41 : _GEN_3112; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3114 = 7'h2a == io_i_rename_table_24 ? io_i_pregs_42 : _GEN_3113; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3115 = 7'h2b == io_i_rename_table_24 ? io_i_pregs_43 : _GEN_3114; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3116 = 7'h2c == io_i_rename_table_24 ? io_i_pregs_44 : _GEN_3115; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3117 = 7'h2d == io_i_rename_table_24 ? io_i_pregs_45 : _GEN_3116; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3118 = 7'h2e == io_i_rename_table_24 ? io_i_pregs_46 : _GEN_3117; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3119 = 7'h2f == io_i_rename_table_24 ? io_i_pregs_47 : _GEN_3118; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3120 = 7'h30 == io_i_rename_table_24 ? io_i_pregs_48 : _GEN_3119; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3121 = 7'h31 == io_i_rename_table_24 ? io_i_pregs_49 : _GEN_3120; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3122 = 7'h32 == io_i_rename_table_24 ? io_i_pregs_50 : _GEN_3121; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3123 = 7'h33 == io_i_rename_table_24 ? io_i_pregs_51 : _GEN_3122; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3124 = 7'h34 == io_i_rename_table_24 ? io_i_pregs_52 : _GEN_3123; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3125 = 7'h35 == io_i_rename_table_24 ? io_i_pregs_53 : _GEN_3124; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3126 = 7'h36 == io_i_rename_table_24 ? io_i_pregs_54 : _GEN_3125; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3127 = 7'h37 == io_i_rename_table_24 ? io_i_pregs_55 : _GEN_3126; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3128 = 7'h38 == io_i_rename_table_24 ? io_i_pregs_56 : _GEN_3127; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3129 = 7'h39 == io_i_rename_table_24 ? io_i_pregs_57 : _GEN_3128; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3130 = 7'h3a == io_i_rename_table_24 ? io_i_pregs_58 : _GEN_3129; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3131 = 7'h3b == io_i_rename_table_24 ? io_i_pregs_59 : _GEN_3130; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3132 = 7'h3c == io_i_rename_table_24 ? io_i_pregs_60 : _GEN_3131; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3133 = 7'h3d == io_i_rename_table_24 ? io_i_pregs_61 : _GEN_3132; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3134 = 7'h3e == io_i_rename_table_24 ? io_i_pregs_62 : _GEN_3133; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3135 = 7'h3f == io_i_rename_table_24 ? io_i_pregs_63 : _GEN_3134; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3136 = 7'h40 == io_i_rename_table_24 ? io_i_pregs_64 : _GEN_3135; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3137 = 7'h41 == io_i_rename_table_24 ? io_i_pregs_65 : _GEN_3136; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3138 = 7'h42 == io_i_rename_table_24 ? io_i_pregs_66 : _GEN_3137; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3139 = 7'h43 == io_i_rename_table_24 ? io_i_pregs_67 : _GEN_3138; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3140 = 7'h44 == io_i_rename_table_24 ? io_i_pregs_68 : _GEN_3139; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3141 = 7'h45 == io_i_rename_table_24 ? io_i_pregs_69 : _GEN_3140; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3142 = 7'h46 == io_i_rename_table_24 ? io_i_pregs_70 : _GEN_3141; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3143 = 7'h47 == io_i_rename_table_24 ? io_i_pregs_71 : _GEN_3142; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3144 = 7'h48 == io_i_rename_table_24 ? io_i_pregs_72 : _GEN_3143; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3145 = 7'h49 == io_i_rename_table_24 ? io_i_pregs_73 : _GEN_3144; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3146 = 7'h4a == io_i_rename_table_24 ? io_i_pregs_74 : _GEN_3145; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3147 = 7'h4b == io_i_rename_table_24 ? io_i_pregs_75 : _GEN_3146; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3148 = 7'h4c == io_i_rename_table_24 ? io_i_pregs_76 : _GEN_3147; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3149 = 7'h4d == io_i_rename_table_24 ? io_i_pregs_77 : _GEN_3148; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3150 = 7'h4e == io_i_rename_table_24 ? io_i_pregs_78 : _GEN_3149; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3151 = 7'h4f == io_i_rename_table_24 ? io_i_pregs_79 : _GEN_3150; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3152 = 7'h50 == io_i_rename_table_24 ? io_i_pregs_80 : _GEN_3151; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3153 = 7'h51 == io_i_rename_table_24 ? io_i_pregs_81 : _GEN_3152; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3154 = 7'h52 == io_i_rename_table_24 ? io_i_pregs_82 : _GEN_3153; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3155 = 7'h53 == io_i_rename_table_24 ? io_i_pregs_83 : _GEN_3154; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3156 = 7'h54 == io_i_rename_table_24 ? io_i_pregs_84 : _GEN_3155; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3157 = 7'h55 == io_i_rename_table_24 ? io_i_pregs_85 : _GEN_3156; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3158 = 7'h56 == io_i_rename_table_24 ? io_i_pregs_86 : _GEN_3157; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3159 = 7'h57 == io_i_rename_table_24 ? io_i_pregs_87 : _GEN_3158; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3160 = 7'h58 == io_i_rename_table_24 ? io_i_pregs_88 : _GEN_3159; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3161 = 7'h59 == io_i_rename_table_24 ? io_i_pregs_89 : _GEN_3160; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3162 = 7'h5a == io_i_rename_table_24 ? io_i_pregs_90 : _GEN_3161; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3163 = 7'h5b == io_i_rename_table_24 ? io_i_pregs_91 : _GEN_3162; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3164 = 7'h5c == io_i_rename_table_24 ? io_i_pregs_92 : _GEN_3163; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3165 = 7'h5d == io_i_rename_table_24 ? io_i_pregs_93 : _GEN_3164; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3166 = 7'h5e == io_i_rename_table_24 ? io_i_pregs_94 : _GEN_3165; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3167 = 7'h5f == io_i_rename_table_24 ? io_i_pregs_95 : _GEN_3166; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3168 = 7'h60 == io_i_rename_table_24 ? io_i_pregs_96 : _GEN_3167; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3169 = 7'h61 == io_i_rename_table_24 ? io_i_pregs_97 : _GEN_3168; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3170 = 7'h62 == io_i_rename_table_24 ? io_i_pregs_98 : _GEN_3169; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3171 = 7'h63 == io_i_rename_table_24 ? io_i_pregs_99 : _GEN_3170; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3172 = 7'h64 == io_i_rename_table_24 ? io_i_pregs_100 : _GEN_3171; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3173 = 7'h65 == io_i_rename_table_24 ? io_i_pregs_101 : _GEN_3172; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3174 = 7'h66 == io_i_rename_table_24 ? io_i_pregs_102 : _GEN_3173; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3175 = 7'h67 == io_i_rename_table_24 ? io_i_pregs_103 : _GEN_3174; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3176 = 7'h68 == io_i_rename_table_24 ? io_i_pregs_104 : _GEN_3175; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3177 = 7'h69 == io_i_rename_table_24 ? io_i_pregs_105 : _GEN_3176; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3178 = 7'h6a == io_i_rename_table_24 ? io_i_pregs_106 : _GEN_3177; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3179 = 7'h6b == io_i_rename_table_24 ? io_i_pregs_107 : _GEN_3178; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3180 = 7'h6c == io_i_rename_table_24 ? io_i_pregs_108 : _GEN_3179; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3181 = 7'h6d == io_i_rename_table_24 ? io_i_pregs_109 : _GEN_3180; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3182 = 7'h6e == io_i_rename_table_24 ? io_i_pregs_110 : _GEN_3181; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3183 = 7'h6f == io_i_rename_table_24 ? io_i_pregs_111 : _GEN_3182; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3184 = 7'h70 == io_i_rename_table_24 ? io_i_pregs_112 : _GEN_3183; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3185 = 7'h71 == io_i_rename_table_24 ? io_i_pregs_113 : _GEN_3184; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3186 = 7'h72 == io_i_rename_table_24 ? io_i_pregs_114 : _GEN_3185; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3187 = 7'h73 == io_i_rename_table_24 ? io_i_pregs_115 : _GEN_3186; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3188 = 7'h74 == io_i_rename_table_24 ? io_i_pregs_116 : _GEN_3187; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3189 = 7'h75 == io_i_rename_table_24 ? io_i_pregs_117 : _GEN_3188; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3190 = 7'h76 == io_i_rename_table_24 ? io_i_pregs_118 : _GEN_3189; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3191 = 7'h77 == io_i_rename_table_24 ? io_i_pregs_119 : _GEN_3190; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3192 = 7'h78 == io_i_rename_table_24 ? io_i_pregs_120 : _GEN_3191; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3193 = 7'h79 == io_i_rename_table_24 ? io_i_pregs_121 : _GEN_3192; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3194 = 7'h7a == io_i_rename_table_24 ? io_i_pregs_122 : _GEN_3193; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3195 = 7'h7b == io_i_rename_table_24 ? io_i_pregs_123 : _GEN_3194; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3196 = 7'h7c == io_i_rename_table_24 ? io_i_pregs_124 : _GEN_3195; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3197 = 7'h7d == io_i_rename_table_24 ? io_i_pregs_125 : _GEN_3196; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3198 = 7'h7e == io_i_rename_table_24 ? io_i_pregs_126 : _GEN_3197; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3201 = 7'h1 == io_i_rename_table_25 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3202 = 7'h2 == io_i_rename_table_25 ? io_i_pregs_2 : _GEN_3201; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3203 = 7'h3 == io_i_rename_table_25 ? io_i_pregs_3 : _GEN_3202; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3204 = 7'h4 == io_i_rename_table_25 ? io_i_pregs_4 : _GEN_3203; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3205 = 7'h5 == io_i_rename_table_25 ? io_i_pregs_5 : _GEN_3204; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3206 = 7'h6 == io_i_rename_table_25 ? io_i_pregs_6 : _GEN_3205; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3207 = 7'h7 == io_i_rename_table_25 ? io_i_pregs_7 : _GEN_3206; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3208 = 7'h8 == io_i_rename_table_25 ? io_i_pregs_8 : _GEN_3207; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3209 = 7'h9 == io_i_rename_table_25 ? io_i_pregs_9 : _GEN_3208; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3210 = 7'ha == io_i_rename_table_25 ? io_i_pregs_10 : _GEN_3209; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3211 = 7'hb == io_i_rename_table_25 ? io_i_pregs_11 : _GEN_3210; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3212 = 7'hc == io_i_rename_table_25 ? io_i_pregs_12 : _GEN_3211; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3213 = 7'hd == io_i_rename_table_25 ? io_i_pregs_13 : _GEN_3212; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3214 = 7'he == io_i_rename_table_25 ? io_i_pregs_14 : _GEN_3213; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3215 = 7'hf == io_i_rename_table_25 ? io_i_pregs_15 : _GEN_3214; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3216 = 7'h10 == io_i_rename_table_25 ? io_i_pregs_16 : _GEN_3215; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3217 = 7'h11 == io_i_rename_table_25 ? io_i_pregs_17 : _GEN_3216; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3218 = 7'h12 == io_i_rename_table_25 ? io_i_pregs_18 : _GEN_3217; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3219 = 7'h13 == io_i_rename_table_25 ? io_i_pregs_19 : _GEN_3218; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3220 = 7'h14 == io_i_rename_table_25 ? io_i_pregs_20 : _GEN_3219; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3221 = 7'h15 == io_i_rename_table_25 ? io_i_pregs_21 : _GEN_3220; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3222 = 7'h16 == io_i_rename_table_25 ? io_i_pregs_22 : _GEN_3221; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3223 = 7'h17 == io_i_rename_table_25 ? io_i_pregs_23 : _GEN_3222; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3224 = 7'h18 == io_i_rename_table_25 ? io_i_pregs_24 : _GEN_3223; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3225 = 7'h19 == io_i_rename_table_25 ? io_i_pregs_25 : _GEN_3224; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3226 = 7'h1a == io_i_rename_table_25 ? io_i_pregs_26 : _GEN_3225; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3227 = 7'h1b == io_i_rename_table_25 ? io_i_pregs_27 : _GEN_3226; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3228 = 7'h1c == io_i_rename_table_25 ? io_i_pregs_28 : _GEN_3227; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3229 = 7'h1d == io_i_rename_table_25 ? io_i_pregs_29 : _GEN_3228; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3230 = 7'h1e == io_i_rename_table_25 ? io_i_pregs_30 : _GEN_3229; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3231 = 7'h1f == io_i_rename_table_25 ? io_i_pregs_31 : _GEN_3230; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3232 = 7'h20 == io_i_rename_table_25 ? io_i_pregs_32 : _GEN_3231; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3233 = 7'h21 == io_i_rename_table_25 ? io_i_pregs_33 : _GEN_3232; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3234 = 7'h22 == io_i_rename_table_25 ? io_i_pregs_34 : _GEN_3233; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3235 = 7'h23 == io_i_rename_table_25 ? io_i_pregs_35 : _GEN_3234; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3236 = 7'h24 == io_i_rename_table_25 ? io_i_pregs_36 : _GEN_3235; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3237 = 7'h25 == io_i_rename_table_25 ? io_i_pregs_37 : _GEN_3236; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3238 = 7'h26 == io_i_rename_table_25 ? io_i_pregs_38 : _GEN_3237; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3239 = 7'h27 == io_i_rename_table_25 ? io_i_pregs_39 : _GEN_3238; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3240 = 7'h28 == io_i_rename_table_25 ? io_i_pregs_40 : _GEN_3239; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3241 = 7'h29 == io_i_rename_table_25 ? io_i_pregs_41 : _GEN_3240; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3242 = 7'h2a == io_i_rename_table_25 ? io_i_pregs_42 : _GEN_3241; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3243 = 7'h2b == io_i_rename_table_25 ? io_i_pregs_43 : _GEN_3242; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3244 = 7'h2c == io_i_rename_table_25 ? io_i_pregs_44 : _GEN_3243; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3245 = 7'h2d == io_i_rename_table_25 ? io_i_pregs_45 : _GEN_3244; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3246 = 7'h2e == io_i_rename_table_25 ? io_i_pregs_46 : _GEN_3245; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3247 = 7'h2f == io_i_rename_table_25 ? io_i_pregs_47 : _GEN_3246; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3248 = 7'h30 == io_i_rename_table_25 ? io_i_pregs_48 : _GEN_3247; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3249 = 7'h31 == io_i_rename_table_25 ? io_i_pregs_49 : _GEN_3248; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3250 = 7'h32 == io_i_rename_table_25 ? io_i_pregs_50 : _GEN_3249; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3251 = 7'h33 == io_i_rename_table_25 ? io_i_pregs_51 : _GEN_3250; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3252 = 7'h34 == io_i_rename_table_25 ? io_i_pregs_52 : _GEN_3251; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3253 = 7'h35 == io_i_rename_table_25 ? io_i_pregs_53 : _GEN_3252; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3254 = 7'h36 == io_i_rename_table_25 ? io_i_pregs_54 : _GEN_3253; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3255 = 7'h37 == io_i_rename_table_25 ? io_i_pregs_55 : _GEN_3254; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3256 = 7'h38 == io_i_rename_table_25 ? io_i_pregs_56 : _GEN_3255; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3257 = 7'h39 == io_i_rename_table_25 ? io_i_pregs_57 : _GEN_3256; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3258 = 7'h3a == io_i_rename_table_25 ? io_i_pregs_58 : _GEN_3257; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3259 = 7'h3b == io_i_rename_table_25 ? io_i_pregs_59 : _GEN_3258; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3260 = 7'h3c == io_i_rename_table_25 ? io_i_pregs_60 : _GEN_3259; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3261 = 7'h3d == io_i_rename_table_25 ? io_i_pregs_61 : _GEN_3260; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3262 = 7'h3e == io_i_rename_table_25 ? io_i_pregs_62 : _GEN_3261; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3263 = 7'h3f == io_i_rename_table_25 ? io_i_pregs_63 : _GEN_3262; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3264 = 7'h40 == io_i_rename_table_25 ? io_i_pregs_64 : _GEN_3263; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3265 = 7'h41 == io_i_rename_table_25 ? io_i_pregs_65 : _GEN_3264; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3266 = 7'h42 == io_i_rename_table_25 ? io_i_pregs_66 : _GEN_3265; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3267 = 7'h43 == io_i_rename_table_25 ? io_i_pregs_67 : _GEN_3266; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3268 = 7'h44 == io_i_rename_table_25 ? io_i_pregs_68 : _GEN_3267; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3269 = 7'h45 == io_i_rename_table_25 ? io_i_pregs_69 : _GEN_3268; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3270 = 7'h46 == io_i_rename_table_25 ? io_i_pregs_70 : _GEN_3269; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3271 = 7'h47 == io_i_rename_table_25 ? io_i_pregs_71 : _GEN_3270; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3272 = 7'h48 == io_i_rename_table_25 ? io_i_pregs_72 : _GEN_3271; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3273 = 7'h49 == io_i_rename_table_25 ? io_i_pregs_73 : _GEN_3272; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3274 = 7'h4a == io_i_rename_table_25 ? io_i_pregs_74 : _GEN_3273; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3275 = 7'h4b == io_i_rename_table_25 ? io_i_pregs_75 : _GEN_3274; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3276 = 7'h4c == io_i_rename_table_25 ? io_i_pregs_76 : _GEN_3275; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3277 = 7'h4d == io_i_rename_table_25 ? io_i_pregs_77 : _GEN_3276; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3278 = 7'h4e == io_i_rename_table_25 ? io_i_pregs_78 : _GEN_3277; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3279 = 7'h4f == io_i_rename_table_25 ? io_i_pregs_79 : _GEN_3278; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3280 = 7'h50 == io_i_rename_table_25 ? io_i_pregs_80 : _GEN_3279; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3281 = 7'h51 == io_i_rename_table_25 ? io_i_pregs_81 : _GEN_3280; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3282 = 7'h52 == io_i_rename_table_25 ? io_i_pregs_82 : _GEN_3281; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3283 = 7'h53 == io_i_rename_table_25 ? io_i_pregs_83 : _GEN_3282; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3284 = 7'h54 == io_i_rename_table_25 ? io_i_pregs_84 : _GEN_3283; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3285 = 7'h55 == io_i_rename_table_25 ? io_i_pregs_85 : _GEN_3284; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3286 = 7'h56 == io_i_rename_table_25 ? io_i_pregs_86 : _GEN_3285; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3287 = 7'h57 == io_i_rename_table_25 ? io_i_pregs_87 : _GEN_3286; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3288 = 7'h58 == io_i_rename_table_25 ? io_i_pregs_88 : _GEN_3287; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3289 = 7'h59 == io_i_rename_table_25 ? io_i_pregs_89 : _GEN_3288; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3290 = 7'h5a == io_i_rename_table_25 ? io_i_pregs_90 : _GEN_3289; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3291 = 7'h5b == io_i_rename_table_25 ? io_i_pregs_91 : _GEN_3290; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3292 = 7'h5c == io_i_rename_table_25 ? io_i_pregs_92 : _GEN_3291; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3293 = 7'h5d == io_i_rename_table_25 ? io_i_pregs_93 : _GEN_3292; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3294 = 7'h5e == io_i_rename_table_25 ? io_i_pregs_94 : _GEN_3293; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3295 = 7'h5f == io_i_rename_table_25 ? io_i_pregs_95 : _GEN_3294; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3296 = 7'h60 == io_i_rename_table_25 ? io_i_pregs_96 : _GEN_3295; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3297 = 7'h61 == io_i_rename_table_25 ? io_i_pregs_97 : _GEN_3296; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3298 = 7'h62 == io_i_rename_table_25 ? io_i_pregs_98 : _GEN_3297; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3299 = 7'h63 == io_i_rename_table_25 ? io_i_pregs_99 : _GEN_3298; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3300 = 7'h64 == io_i_rename_table_25 ? io_i_pregs_100 : _GEN_3299; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3301 = 7'h65 == io_i_rename_table_25 ? io_i_pregs_101 : _GEN_3300; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3302 = 7'h66 == io_i_rename_table_25 ? io_i_pregs_102 : _GEN_3301; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3303 = 7'h67 == io_i_rename_table_25 ? io_i_pregs_103 : _GEN_3302; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3304 = 7'h68 == io_i_rename_table_25 ? io_i_pregs_104 : _GEN_3303; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3305 = 7'h69 == io_i_rename_table_25 ? io_i_pregs_105 : _GEN_3304; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3306 = 7'h6a == io_i_rename_table_25 ? io_i_pregs_106 : _GEN_3305; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3307 = 7'h6b == io_i_rename_table_25 ? io_i_pregs_107 : _GEN_3306; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3308 = 7'h6c == io_i_rename_table_25 ? io_i_pregs_108 : _GEN_3307; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3309 = 7'h6d == io_i_rename_table_25 ? io_i_pregs_109 : _GEN_3308; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3310 = 7'h6e == io_i_rename_table_25 ? io_i_pregs_110 : _GEN_3309; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3311 = 7'h6f == io_i_rename_table_25 ? io_i_pregs_111 : _GEN_3310; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3312 = 7'h70 == io_i_rename_table_25 ? io_i_pregs_112 : _GEN_3311; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3313 = 7'h71 == io_i_rename_table_25 ? io_i_pregs_113 : _GEN_3312; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3314 = 7'h72 == io_i_rename_table_25 ? io_i_pregs_114 : _GEN_3313; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3315 = 7'h73 == io_i_rename_table_25 ? io_i_pregs_115 : _GEN_3314; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3316 = 7'h74 == io_i_rename_table_25 ? io_i_pregs_116 : _GEN_3315; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3317 = 7'h75 == io_i_rename_table_25 ? io_i_pregs_117 : _GEN_3316; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3318 = 7'h76 == io_i_rename_table_25 ? io_i_pregs_118 : _GEN_3317; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3319 = 7'h77 == io_i_rename_table_25 ? io_i_pregs_119 : _GEN_3318; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3320 = 7'h78 == io_i_rename_table_25 ? io_i_pregs_120 : _GEN_3319; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3321 = 7'h79 == io_i_rename_table_25 ? io_i_pregs_121 : _GEN_3320; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3322 = 7'h7a == io_i_rename_table_25 ? io_i_pregs_122 : _GEN_3321; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3323 = 7'h7b == io_i_rename_table_25 ? io_i_pregs_123 : _GEN_3322; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3324 = 7'h7c == io_i_rename_table_25 ? io_i_pregs_124 : _GEN_3323; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3325 = 7'h7d == io_i_rename_table_25 ? io_i_pregs_125 : _GEN_3324; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3326 = 7'h7e == io_i_rename_table_25 ? io_i_pregs_126 : _GEN_3325; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3329 = 7'h1 == io_i_rename_table_26 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3330 = 7'h2 == io_i_rename_table_26 ? io_i_pregs_2 : _GEN_3329; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3331 = 7'h3 == io_i_rename_table_26 ? io_i_pregs_3 : _GEN_3330; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3332 = 7'h4 == io_i_rename_table_26 ? io_i_pregs_4 : _GEN_3331; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3333 = 7'h5 == io_i_rename_table_26 ? io_i_pregs_5 : _GEN_3332; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3334 = 7'h6 == io_i_rename_table_26 ? io_i_pregs_6 : _GEN_3333; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3335 = 7'h7 == io_i_rename_table_26 ? io_i_pregs_7 : _GEN_3334; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3336 = 7'h8 == io_i_rename_table_26 ? io_i_pregs_8 : _GEN_3335; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3337 = 7'h9 == io_i_rename_table_26 ? io_i_pregs_9 : _GEN_3336; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3338 = 7'ha == io_i_rename_table_26 ? io_i_pregs_10 : _GEN_3337; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3339 = 7'hb == io_i_rename_table_26 ? io_i_pregs_11 : _GEN_3338; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3340 = 7'hc == io_i_rename_table_26 ? io_i_pregs_12 : _GEN_3339; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3341 = 7'hd == io_i_rename_table_26 ? io_i_pregs_13 : _GEN_3340; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3342 = 7'he == io_i_rename_table_26 ? io_i_pregs_14 : _GEN_3341; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3343 = 7'hf == io_i_rename_table_26 ? io_i_pregs_15 : _GEN_3342; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3344 = 7'h10 == io_i_rename_table_26 ? io_i_pregs_16 : _GEN_3343; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3345 = 7'h11 == io_i_rename_table_26 ? io_i_pregs_17 : _GEN_3344; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3346 = 7'h12 == io_i_rename_table_26 ? io_i_pregs_18 : _GEN_3345; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3347 = 7'h13 == io_i_rename_table_26 ? io_i_pregs_19 : _GEN_3346; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3348 = 7'h14 == io_i_rename_table_26 ? io_i_pregs_20 : _GEN_3347; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3349 = 7'h15 == io_i_rename_table_26 ? io_i_pregs_21 : _GEN_3348; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3350 = 7'h16 == io_i_rename_table_26 ? io_i_pregs_22 : _GEN_3349; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3351 = 7'h17 == io_i_rename_table_26 ? io_i_pregs_23 : _GEN_3350; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3352 = 7'h18 == io_i_rename_table_26 ? io_i_pregs_24 : _GEN_3351; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3353 = 7'h19 == io_i_rename_table_26 ? io_i_pregs_25 : _GEN_3352; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3354 = 7'h1a == io_i_rename_table_26 ? io_i_pregs_26 : _GEN_3353; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3355 = 7'h1b == io_i_rename_table_26 ? io_i_pregs_27 : _GEN_3354; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3356 = 7'h1c == io_i_rename_table_26 ? io_i_pregs_28 : _GEN_3355; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3357 = 7'h1d == io_i_rename_table_26 ? io_i_pregs_29 : _GEN_3356; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3358 = 7'h1e == io_i_rename_table_26 ? io_i_pregs_30 : _GEN_3357; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3359 = 7'h1f == io_i_rename_table_26 ? io_i_pregs_31 : _GEN_3358; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3360 = 7'h20 == io_i_rename_table_26 ? io_i_pregs_32 : _GEN_3359; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3361 = 7'h21 == io_i_rename_table_26 ? io_i_pregs_33 : _GEN_3360; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3362 = 7'h22 == io_i_rename_table_26 ? io_i_pregs_34 : _GEN_3361; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3363 = 7'h23 == io_i_rename_table_26 ? io_i_pregs_35 : _GEN_3362; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3364 = 7'h24 == io_i_rename_table_26 ? io_i_pregs_36 : _GEN_3363; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3365 = 7'h25 == io_i_rename_table_26 ? io_i_pregs_37 : _GEN_3364; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3366 = 7'h26 == io_i_rename_table_26 ? io_i_pregs_38 : _GEN_3365; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3367 = 7'h27 == io_i_rename_table_26 ? io_i_pregs_39 : _GEN_3366; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3368 = 7'h28 == io_i_rename_table_26 ? io_i_pregs_40 : _GEN_3367; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3369 = 7'h29 == io_i_rename_table_26 ? io_i_pregs_41 : _GEN_3368; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3370 = 7'h2a == io_i_rename_table_26 ? io_i_pregs_42 : _GEN_3369; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3371 = 7'h2b == io_i_rename_table_26 ? io_i_pregs_43 : _GEN_3370; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3372 = 7'h2c == io_i_rename_table_26 ? io_i_pregs_44 : _GEN_3371; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3373 = 7'h2d == io_i_rename_table_26 ? io_i_pregs_45 : _GEN_3372; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3374 = 7'h2e == io_i_rename_table_26 ? io_i_pregs_46 : _GEN_3373; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3375 = 7'h2f == io_i_rename_table_26 ? io_i_pregs_47 : _GEN_3374; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3376 = 7'h30 == io_i_rename_table_26 ? io_i_pregs_48 : _GEN_3375; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3377 = 7'h31 == io_i_rename_table_26 ? io_i_pregs_49 : _GEN_3376; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3378 = 7'h32 == io_i_rename_table_26 ? io_i_pregs_50 : _GEN_3377; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3379 = 7'h33 == io_i_rename_table_26 ? io_i_pregs_51 : _GEN_3378; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3380 = 7'h34 == io_i_rename_table_26 ? io_i_pregs_52 : _GEN_3379; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3381 = 7'h35 == io_i_rename_table_26 ? io_i_pregs_53 : _GEN_3380; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3382 = 7'h36 == io_i_rename_table_26 ? io_i_pregs_54 : _GEN_3381; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3383 = 7'h37 == io_i_rename_table_26 ? io_i_pregs_55 : _GEN_3382; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3384 = 7'h38 == io_i_rename_table_26 ? io_i_pregs_56 : _GEN_3383; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3385 = 7'h39 == io_i_rename_table_26 ? io_i_pregs_57 : _GEN_3384; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3386 = 7'h3a == io_i_rename_table_26 ? io_i_pregs_58 : _GEN_3385; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3387 = 7'h3b == io_i_rename_table_26 ? io_i_pregs_59 : _GEN_3386; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3388 = 7'h3c == io_i_rename_table_26 ? io_i_pregs_60 : _GEN_3387; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3389 = 7'h3d == io_i_rename_table_26 ? io_i_pregs_61 : _GEN_3388; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3390 = 7'h3e == io_i_rename_table_26 ? io_i_pregs_62 : _GEN_3389; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3391 = 7'h3f == io_i_rename_table_26 ? io_i_pregs_63 : _GEN_3390; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3392 = 7'h40 == io_i_rename_table_26 ? io_i_pregs_64 : _GEN_3391; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3393 = 7'h41 == io_i_rename_table_26 ? io_i_pregs_65 : _GEN_3392; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3394 = 7'h42 == io_i_rename_table_26 ? io_i_pregs_66 : _GEN_3393; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3395 = 7'h43 == io_i_rename_table_26 ? io_i_pregs_67 : _GEN_3394; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3396 = 7'h44 == io_i_rename_table_26 ? io_i_pregs_68 : _GEN_3395; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3397 = 7'h45 == io_i_rename_table_26 ? io_i_pregs_69 : _GEN_3396; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3398 = 7'h46 == io_i_rename_table_26 ? io_i_pregs_70 : _GEN_3397; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3399 = 7'h47 == io_i_rename_table_26 ? io_i_pregs_71 : _GEN_3398; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3400 = 7'h48 == io_i_rename_table_26 ? io_i_pregs_72 : _GEN_3399; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3401 = 7'h49 == io_i_rename_table_26 ? io_i_pregs_73 : _GEN_3400; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3402 = 7'h4a == io_i_rename_table_26 ? io_i_pregs_74 : _GEN_3401; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3403 = 7'h4b == io_i_rename_table_26 ? io_i_pregs_75 : _GEN_3402; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3404 = 7'h4c == io_i_rename_table_26 ? io_i_pregs_76 : _GEN_3403; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3405 = 7'h4d == io_i_rename_table_26 ? io_i_pregs_77 : _GEN_3404; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3406 = 7'h4e == io_i_rename_table_26 ? io_i_pregs_78 : _GEN_3405; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3407 = 7'h4f == io_i_rename_table_26 ? io_i_pregs_79 : _GEN_3406; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3408 = 7'h50 == io_i_rename_table_26 ? io_i_pregs_80 : _GEN_3407; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3409 = 7'h51 == io_i_rename_table_26 ? io_i_pregs_81 : _GEN_3408; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3410 = 7'h52 == io_i_rename_table_26 ? io_i_pregs_82 : _GEN_3409; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3411 = 7'h53 == io_i_rename_table_26 ? io_i_pregs_83 : _GEN_3410; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3412 = 7'h54 == io_i_rename_table_26 ? io_i_pregs_84 : _GEN_3411; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3413 = 7'h55 == io_i_rename_table_26 ? io_i_pregs_85 : _GEN_3412; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3414 = 7'h56 == io_i_rename_table_26 ? io_i_pregs_86 : _GEN_3413; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3415 = 7'h57 == io_i_rename_table_26 ? io_i_pregs_87 : _GEN_3414; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3416 = 7'h58 == io_i_rename_table_26 ? io_i_pregs_88 : _GEN_3415; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3417 = 7'h59 == io_i_rename_table_26 ? io_i_pregs_89 : _GEN_3416; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3418 = 7'h5a == io_i_rename_table_26 ? io_i_pregs_90 : _GEN_3417; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3419 = 7'h5b == io_i_rename_table_26 ? io_i_pregs_91 : _GEN_3418; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3420 = 7'h5c == io_i_rename_table_26 ? io_i_pregs_92 : _GEN_3419; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3421 = 7'h5d == io_i_rename_table_26 ? io_i_pregs_93 : _GEN_3420; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3422 = 7'h5e == io_i_rename_table_26 ? io_i_pregs_94 : _GEN_3421; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3423 = 7'h5f == io_i_rename_table_26 ? io_i_pregs_95 : _GEN_3422; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3424 = 7'h60 == io_i_rename_table_26 ? io_i_pregs_96 : _GEN_3423; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3425 = 7'h61 == io_i_rename_table_26 ? io_i_pregs_97 : _GEN_3424; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3426 = 7'h62 == io_i_rename_table_26 ? io_i_pregs_98 : _GEN_3425; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3427 = 7'h63 == io_i_rename_table_26 ? io_i_pregs_99 : _GEN_3426; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3428 = 7'h64 == io_i_rename_table_26 ? io_i_pregs_100 : _GEN_3427; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3429 = 7'h65 == io_i_rename_table_26 ? io_i_pregs_101 : _GEN_3428; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3430 = 7'h66 == io_i_rename_table_26 ? io_i_pregs_102 : _GEN_3429; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3431 = 7'h67 == io_i_rename_table_26 ? io_i_pregs_103 : _GEN_3430; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3432 = 7'h68 == io_i_rename_table_26 ? io_i_pregs_104 : _GEN_3431; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3433 = 7'h69 == io_i_rename_table_26 ? io_i_pregs_105 : _GEN_3432; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3434 = 7'h6a == io_i_rename_table_26 ? io_i_pregs_106 : _GEN_3433; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3435 = 7'h6b == io_i_rename_table_26 ? io_i_pregs_107 : _GEN_3434; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3436 = 7'h6c == io_i_rename_table_26 ? io_i_pregs_108 : _GEN_3435; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3437 = 7'h6d == io_i_rename_table_26 ? io_i_pregs_109 : _GEN_3436; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3438 = 7'h6e == io_i_rename_table_26 ? io_i_pregs_110 : _GEN_3437; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3439 = 7'h6f == io_i_rename_table_26 ? io_i_pregs_111 : _GEN_3438; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3440 = 7'h70 == io_i_rename_table_26 ? io_i_pregs_112 : _GEN_3439; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3441 = 7'h71 == io_i_rename_table_26 ? io_i_pregs_113 : _GEN_3440; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3442 = 7'h72 == io_i_rename_table_26 ? io_i_pregs_114 : _GEN_3441; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3443 = 7'h73 == io_i_rename_table_26 ? io_i_pregs_115 : _GEN_3442; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3444 = 7'h74 == io_i_rename_table_26 ? io_i_pregs_116 : _GEN_3443; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3445 = 7'h75 == io_i_rename_table_26 ? io_i_pregs_117 : _GEN_3444; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3446 = 7'h76 == io_i_rename_table_26 ? io_i_pregs_118 : _GEN_3445; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3447 = 7'h77 == io_i_rename_table_26 ? io_i_pregs_119 : _GEN_3446; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3448 = 7'h78 == io_i_rename_table_26 ? io_i_pregs_120 : _GEN_3447; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3449 = 7'h79 == io_i_rename_table_26 ? io_i_pregs_121 : _GEN_3448; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3450 = 7'h7a == io_i_rename_table_26 ? io_i_pregs_122 : _GEN_3449; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3451 = 7'h7b == io_i_rename_table_26 ? io_i_pregs_123 : _GEN_3450; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3452 = 7'h7c == io_i_rename_table_26 ? io_i_pregs_124 : _GEN_3451; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3453 = 7'h7d == io_i_rename_table_26 ? io_i_pregs_125 : _GEN_3452; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3454 = 7'h7e == io_i_rename_table_26 ? io_i_pregs_126 : _GEN_3453; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3457 = 7'h1 == io_i_rename_table_27 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3458 = 7'h2 == io_i_rename_table_27 ? io_i_pregs_2 : _GEN_3457; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3459 = 7'h3 == io_i_rename_table_27 ? io_i_pregs_3 : _GEN_3458; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3460 = 7'h4 == io_i_rename_table_27 ? io_i_pregs_4 : _GEN_3459; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3461 = 7'h5 == io_i_rename_table_27 ? io_i_pregs_5 : _GEN_3460; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3462 = 7'h6 == io_i_rename_table_27 ? io_i_pregs_6 : _GEN_3461; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3463 = 7'h7 == io_i_rename_table_27 ? io_i_pregs_7 : _GEN_3462; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3464 = 7'h8 == io_i_rename_table_27 ? io_i_pregs_8 : _GEN_3463; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3465 = 7'h9 == io_i_rename_table_27 ? io_i_pregs_9 : _GEN_3464; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3466 = 7'ha == io_i_rename_table_27 ? io_i_pregs_10 : _GEN_3465; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3467 = 7'hb == io_i_rename_table_27 ? io_i_pregs_11 : _GEN_3466; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3468 = 7'hc == io_i_rename_table_27 ? io_i_pregs_12 : _GEN_3467; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3469 = 7'hd == io_i_rename_table_27 ? io_i_pregs_13 : _GEN_3468; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3470 = 7'he == io_i_rename_table_27 ? io_i_pregs_14 : _GEN_3469; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3471 = 7'hf == io_i_rename_table_27 ? io_i_pregs_15 : _GEN_3470; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3472 = 7'h10 == io_i_rename_table_27 ? io_i_pregs_16 : _GEN_3471; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3473 = 7'h11 == io_i_rename_table_27 ? io_i_pregs_17 : _GEN_3472; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3474 = 7'h12 == io_i_rename_table_27 ? io_i_pregs_18 : _GEN_3473; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3475 = 7'h13 == io_i_rename_table_27 ? io_i_pregs_19 : _GEN_3474; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3476 = 7'h14 == io_i_rename_table_27 ? io_i_pregs_20 : _GEN_3475; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3477 = 7'h15 == io_i_rename_table_27 ? io_i_pregs_21 : _GEN_3476; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3478 = 7'h16 == io_i_rename_table_27 ? io_i_pregs_22 : _GEN_3477; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3479 = 7'h17 == io_i_rename_table_27 ? io_i_pregs_23 : _GEN_3478; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3480 = 7'h18 == io_i_rename_table_27 ? io_i_pregs_24 : _GEN_3479; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3481 = 7'h19 == io_i_rename_table_27 ? io_i_pregs_25 : _GEN_3480; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3482 = 7'h1a == io_i_rename_table_27 ? io_i_pregs_26 : _GEN_3481; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3483 = 7'h1b == io_i_rename_table_27 ? io_i_pregs_27 : _GEN_3482; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3484 = 7'h1c == io_i_rename_table_27 ? io_i_pregs_28 : _GEN_3483; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3485 = 7'h1d == io_i_rename_table_27 ? io_i_pregs_29 : _GEN_3484; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3486 = 7'h1e == io_i_rename_table_27 ? io_i_pregs_30 : _GEN_3485; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3487 = 7'h1f == io_i_rename_table_27 ? io_i_pregs_31 : _GEN_3486; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3488 = 7'h20 == io_i_rename_table_27 ? io_i_pregs_32 : _GEN_3487; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3489 = 7'h21 == io_i_rename_table_27 ? io_i_pregs_33 : _GEN_3488; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3490 = 7'h22 == io_i_rename_table_27 ? io_i_pregs_34 : _GEN_3489; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3491 = 7'h23 == io_i_rename_table_27 ? io_i_pregs_35 : _GEN_3490; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3492 = 7'h24 == io_i_rename_table_27 ? io_i_pregs_36 : _GEN_3491; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3493 = 7'h25 == io_i_rename_table_27 ? io_i_pregs_37 : _GEN_3492; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3494 = 7'h26 == io_i_rename_table_27 ? io_i_pregs_38 : _GEN_3493; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3495 = 7'h27 == io_i_rename_table_27 ? io_i_pregs_39 : _GEN_3494; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3496 = 7'h28 == io_i_rename_table_27 ? io_i_pregs_40 : _GEN_3495; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3497 = 7'h29 == io_i_rename_table_27 ? io_i_pregs_41 : _GEN_3496; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3498 = 7'h2a == io_i_rename_table_27 ? io_i_pregs_42 : _GEN_3497; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3499 = 7'h2b == io_i_rename_table_27 ? io_i_pregs_43 : _GEN_3498; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3500 = 7'h2c == io_i_rename_table_27 ? io_i_pregs_44 : _GEN_3499; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3501 = 7'h2d == io_i_rename_table_27 ? io_i_pregs_45 : _GEN_3500; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3502 = 7'h2e == io_i_rename_table_27 ? io_i_pregs_46 : _GEN_3501; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3503 = 7'h2f == io_i_rename_table_27 ? io_i_pregs_47 : _GEN_3502; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3504 = 7'h30 == io_i_rename_table_27 ? io_i_pregs_48 : _GEN_3503; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3505 = 7'h31 == io_i_rename_table_27 ? io_i_pregs_49 : _GEN_3504; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3506 = 7'h32 == io_i_rename_table_27 ? io_i_pregs_50 : _GEN_3505; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3507 = 7'h33 == io_i_rename_table_27 ? io_i_pregs_51 : _GEN_3506; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3508 = 7'h34 == io_i_rename_table_27 ? io_i_pregs_52 : _GEN_3507; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3509 = 7'h35 == io_i_rename_table_27 ? io_i_pregs_53 : _GEN_3508; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3510 = 7'h36 == io_i_rename_table_27 ? io_i_pregs_54 : _GEN_3509; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3511 = 7'h37 == io_i_rename_table_27 ? io_i_pregs_55 : _GEN_3510; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3512 = 7'h38 == io_i_rename_table_27 ? io_i_pregs_56 : _GEN_3511; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3513 = 7'h39 == io_i_rename_table_27 ? io_i_pregs_57 : _GEN_3512; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3514 = 7'h3a == io_i_rename_table_27 ? io_i_pregs_58 : _GEN_3513; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3515 = 7'h3b == io_i_rename_table_27 ? io_i_pregs_59 : _GEN_3514; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3516 = 7'h3c == io_i_rename_table_27 ? io_i_pregs_60 : _GEN_3515; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3517 = 7'h3d == io_i_rename_table_27 ? io_i_pregs_61 : _GEN_3516; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3518 = 7'h3e == io_i_rename_table_27 ? io_i_pregs_62 : _GEN_3517; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3519 = 7'h3f == io_i_rename_table_27 ? io_i_pregs_63 : _GEN_3518; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3520 = 7'h40 == io_i_rename_table_27 ? io_i_pregs_64 : _GEN_3519; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3521 = 7'h41 == io_i_rename_table_27 ? io_i_pregs_65 : _GEN_3520; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3522 = 7'h42 == io_i_rename_table_27 ? io_i_pregs_66 : _GEN_3521; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3523 = 7'h43 == io_i_rename_table_27 ? io_i_pregs_67 : _GEN_3522; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3524 = 7'h44 == io_i_rename_table_27 ? io_i_pregs_68 : _GEN_3523; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3525 = 7'h45 == io_i_rename_table_27 ? io_i_pregs_69 : _GEN_3524; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3526 = 7'h46 == io_i_rename_table_27 ? io_i_pregs_70 : _GEN_3525; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3527 = 7'h47 == io_i_rename_table_27 ? io_i_pregs_71 : _GEN_3526; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3528 = 7'h48 == io_i_rename_table_27 ? io_i_pregs_72 : _GEN_3527; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3529 = 7'h49 == io_i_rename_table_27 ? io_i_pregs_73 : _GEN_3528; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3530 = 7'h4a == io_i_rename_table_27 ? io_i_pregs_74 : _GEN_3529; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3531 = 7'h4b == io_i_rename_table_27 ? io_i_pregs_75 : _GEN_3530; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3532 = 7'h4c == io_i_rename_table_27 ? io_i_pregs_76 : _GEN_3531; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3533 = 7'h4d == io_i_rename_table_27 ? io_i_pregs_77 : _GEN_3532; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3534 = 7'h4e == io_i_rename_table_27 ? io_i_pregs_78 : _GEN_3533; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3535 = 7'h4f == io_i_rename_table_27 ? io_i_pregs_79 : _GEN_3534; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3536 = 7'h50 == io_i_rename_table_27 ? io_i_pregs_80 : _GEN_3535; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3537 = 7'h51 == io_i_rename_table_27 ? io_i_pregs_81 : _GEN_3536; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3538 = 7'h52 == io_i_rename_table_27 ? io_i_pregs_82 : _GEN_3537; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3539 = 7'h53 == io_i_rename_table_27 ? io_i_pregs_83 : _GEN_3538; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3540 = 7'h54 == io_i_rename_table_27 ? io_i_pregs_84 : _GEN_3539; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3541 = 7'h55 == io_i_rename_table_27 ? io_i_pregs_85 : _GEN_3540; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3542 = 7'h56 == io_i_rename_table_27 ? io_i_pregs_86 : _GEN_3541; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3543 = 7'h57 == io_i_rename_table_27 ? io_i_pregs_87 : _GEN_3542; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3544 = 7'h58 == io_i_rename_table_27 ? io_i_pregs_88 : _GEN_3543; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3545 = 7'h59 == io_i_rename_table_27 ? io_i_pregs_89 : _GEN_3544; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3546 = 7'h5a == io_i_rename_table_27 ? io_i_pregs_90 : _GEN_3545; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3547 = 7'h5b == io_i_rename_table_27 ? io_i_pregs_91 : _GEN_3546; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3548 = 7'h5c == io_i_rename_table_27 ? io_i_pregs_92 : _GEN_3547; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3549 = 7'h5d == io_i_rename_table_27 ? io_i_pregs_93 : _GEN_3548; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3550 = 7'h5e == io_i_rename_table_27 ? io_i_pregs_94 : _GEN_3549; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3551 = 7'h5f == io_i_rename_table_27 ? io_i_pregs_95 : _GEN_3550; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3552 = 7'h60 == io_i_rename_table_27 ? io_i_pregs_96 : _GEN_3551; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3553 = 7'h61 == io_i_rename_table_27 ? io_i_pregs_97 : _GEN_3552; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3554 = 7'h62 == io_i_rename_table_27 ? io_i_pregs_98 : _GEN_3553; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3555 = 7'h63 == io_i_rename_table_27 ? io_i_pregs_99 : _GEN_3554; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3556 = 7'h64 == io_i_rename_table_27 ? io_i_pregs_100 : _GEN_3555; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3557 = 7'h65 == io_i_rename_table_27 ? io_i_pregs_101 : _GEN_3556; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3558 = 7'h66 == io_i_rename_table_27 ? io_i_pregs_102 : _GEN_3557; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3559 = 7'h67 == io_i_rename_table_27 ? io_i_pregs_103 : _GEN_3558; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3560 = 7'h68 == io_i_rename_table_27 ? io_i_pregs_104 : _GEN_3559; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3561 = 7'h69 == io_i_rename_table_27 ? io_i_pregs_105 : _GEN_3560; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3562 = 7'h6a == io_i_rename_table_27 ? io_i_pregs_106 : _GEN_3561; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3563 = 7'h6b == io_i_rename_table_27 ? io_i_pregs_107 : _GEN_3562; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3564 = 7'h6c == io_i_rename_table_27 ? io_i_pregs_108 : _GEN_3563; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3565 = 7'h6d == io_i_rename_table_27 ? io_i_pregs_109 : _GEN_3564; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3566 = 7'h6e == io_i_rename_table_27 ? io_i_pregs_110 : _GEN_3565; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3567 = 7'h6f == io_i_rename_table_27 ? io_i_pregs_111 : _GEN_3566; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3568 = 7'h70 == io_i_rename_table_27 ? io_i_pregs_112 : _GEN_3567; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3569 = 7'h71 == io_i_rename_table_27 ? io_i_pregs_113 : _GEN_3568; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3570 = 7'h72 == io_i_rename_table_27 ? io_i_pregs_114 : _GEN_3569; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3571 = 7'h73 == io_i_rename_table_27 ? io_i_pregs_115 : _GEN_3570; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3572 = 7'h74 == io_i_rename_table_27 ? io_i_pregs_116 : _GEN_3571; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3573 = 7'h75 == io_i_rename_table_27 ? io_i_pregs_117 : _GEN_3572; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3574 = 7'h76 == io_i_rename_table_27 ? io_i_pregs_118 : _GEN_3573; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3575 = 7'h77 == io_i_rename_table_27 ? io_i_pregs_119 : _GEN_3574; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3576 = 7'h78 == io_i_rename_table_27 ? io_i_pregs_120 : _GEN_3575; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3577 = 7'h79 == io_i_rename_table_27 ? io_i_pregs_121 : _GEN_3576; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3578 = 7'h7a == io_i_rename_table_27 ? io_i_pregs_122 : _GEN_3577; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3579 = 7'h7b == io_i_rename_table_27 ? io_i_pregs_123 : _GEN_3578; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3580 = 7'h7c == io_i_rename_table_27 ? io_i_pregs_124 : _GEN_3579; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3581 = 7'h7d == io_i_rename_table_27 ? io_i_pregs_125 : _GEN_3580; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3582 = 7'h7e == io_i_rename_table_27 ? io_i_pregs_126 : _GEN_3581; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3585 = 7'h1 == io_i_rename_table_28 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3586 = 7'h2 == io_i_rename_table_28 ? io_i_pregs_2 : _GEN_3585; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3587 = 7'h3 == io_i_rename_table_28 ? io_i_pregs_3 : _GEN_3586; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3588 = 7'h4 == io_i_rename_table_28 ? io_i_pregs_4 : _GEN_3587; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3589 = 7'h5 == io_i_rename_table_28 ? io_i_pregs_5 : _GEN_3588; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3590 = 7'h6 == io_i_rename_table_28 ? io_i_pregs_6 : _GEN_3589; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3591 = 7'h7 == io_i_rename_table_28 ? io_i_pregs_7 : _GEN_3590; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3592 = 7'h8 == io_i_rename_table_28 ? io_i_pregs_8 : _GEN_3591; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3593 = 7'h9 == io_i_rename_table_28 ? io_i_pregs_9 : _GEN_3592; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3594 = 7'ha == io_i_rename_table_28 ? io_i_pregs_10 : _GEN_3593; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3595 = 7'hb == io_i_rename_table_28 ? io_i_pregs_11 : _GEN_3594; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3596 = 7'hc == io_i_rename_table_28 ? io_i_pregs_12 : _GEN_3595; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3597 = 7'hd == io_i_rename_table_28 ? io_i_pregs_13 : _GEN_3596; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3598 = 7'he == io_i_rename_table_28 ? io_i_pregs_14 : _GEN_3597; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3599 = 7'hf == io_i_rename_table_28 ? io_i_pregs_15 : _GEN_3598; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3600 = 7'h10 == io_i_rename_table_28 ? io_i_pregs_16 : _GEN_3599; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3601 = 7'h11 == io_i_rename_table_28 ? io_i_pregs_17 : _GEN_3600; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3602 = 7'h12 == io_i_rename_table_28 ? io_i_pregs_18 : _GEN_3601; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3603 = 7'h13 == io_i_rename_table_28 ? io_i_pregs_19 : _GEN_3602; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3604 = 7'h14 == io_i_rename_table_28 ? io_i_pregs_20 : _GEN_3603; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3605 = 7'h15 == io_i_rename_table_28 ? io_i_pregs_21 : _GEN_3604; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3606 = 7'h16 == io_i_rename_table_28 ? io_i_pregs_22 : _GEN_3605; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3607 = 7'h17 == io_i_rename_table_28 ? io_i_pregs_23 : _GEN_3606; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3608 = 7'h18 == io_i_rename_table_28 ? io_i_pregs_24 : _GEN_3607; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3609 = 7'h19 == io_i_rename_table_28 ? io_i_pregs_25 : _GEN_3608; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3610 = 7'h1a == io_i_rename_table_28 ? io_i_pregs_26 : _GEN_3609; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3611 = 7'h1b == io_i_rename_table_28 ? io_i_pregs_27 : _GEN_3610; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3612 = 7'h1c == io_i_rename_table_28 ? io_i_pregs_28 : _GEN_3611; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3613 = 7'h1d == io_i_rename_table_28 ? io_i_pregs_29 : _GEN_3612; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3614 = 7'h1e == io_i_rename_table_28 ? io_i_pregs_30 : _GEN_3613; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3615 = 7'h1f == io_i_rename_table_28 ? io_i_pregs_31 : _GEN_3614; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3616 = 7'h20 == io_i_rename_table_28 ? io_i_pregs_32 : _GEN_3615; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3617 = 7'h21 == io_i_rename_table_28 ? io_i_pregs_33 : _GEN_3616; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3618 = 7'h22 == io_i_rename_table_28 ? io_i_pregs_34 : _GEN_3617; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3619 = 7'h23 == io_i_rename_table_28 ? io_i_pregs_35 : _GEN_3618; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3620 = 7'h24 == io_i_rename_table_28 ? io_i_pregs_36 : _GEN_3619; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3621 = 7'h25 == io_i_rename_table_28 ? io_i_pregs_37 : _GEN_3620; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3622 = 7'h26 == io_i_rename_table_28 ? io_i_pregs_38 : _GEN_3621; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3623 = 7'h27 == io_i_rename_table_28 ? io_i_pregs_39 : _GEN_3622; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3624 = 7'h28 == io_i_rename_table_28 ? io_i_pregs_40 : _GEN_3623; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3625 = 7'h29 == io_i_rename_table_28 ? io_i_pregs_41 : _GEN_3624; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3626 = 7'h2a == io_i_rename_table_28 ? io_i_pregs_42 : _GEN_3625; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3627 = 7'h2b == io_i_rename_table_28 ? io_i_pregs_43 : _GEN_3626; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3628 = 7'h2c == io_i_rename_table_28 ? io_i_pregs_44 : _GEN_3627; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3629 = 7'h2d == io_i_rename_table_28 ? io_i_pregs_45 : _GEN_3628; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3630 = 7'h2e == io_i_rename_table_28 ? io_i_pregs_46 : _GEN_3629; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3631 = 7'h2f == io_i_rename_table_28 ? io_i_pregs_47 : _GEN_3630; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3632 = 7'h30 == io_i_rename_table_28 ? io_i_pregs_48 : _GEN_3631; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3633 = 7'h31 == io_i_rename_table_28 ? io_i_pregs_49 : _GEN_3632; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3634 = 7'h32 == io_i_rename_table_28 ? io_i_pregs_50 : _GEN_3633; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3635 = 7'h33 == io_i_rename_table_28 ? io_i_pregs_51 : _GEN_3634; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3636 = 7'h34 == io_i_rename_table_28 ? io_i_pregs_52 : _GEN_3635; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3637 = 7'h35 == io_i_rename_table_28 ? io_i_pregs_53 : _GEN_3636; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3638 = 7'h36 == io_i_rename_table_28 ? io_i_pregs_54 : _GEN_3637; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3639 = 7'h37 == io_i_rename_table_28 ? io_i_pregs_55 : _GEN_3638; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3640 = 7'h38 == io_i_rename_table_28 ? io_i_pregs_56 : _GEN_3639; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3641 = 7'h39 == io_i_rename_table_28 ? io_i_pregs_57 : _GEN_3640; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3642 = 7'h3a == io_i_rename_table_28 ? io_i_pregs_58 : _GEN_3641; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3643 = 7'h3b == io_i_rename_table_28 ? io_i_pregs_59 : _GEN_3642; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3644 = 7'h3c == io_i_rename_table_28 ? io_i_pregs_60 : _GEN_3643; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3645 = 7'h3d == io_i_rename_table_28 ? io_i_pregs_61 : _GEN_3644; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3646 = 7'h3e == io_i_rename_table_28 ? io_i_pregs_62 : _GEN_3645; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3647 = 7'h3f == io_i_rename_table_28 ? io_i_pregs_63 : _GEN_3646; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3648 = 7'h40 == io_i_rename_table_28 ? io_i_pregs_64 : _GEN_3647; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3649 = 7'h41 == io_i_rename_table_28 ? io_i_pregs_65 : _GEN_3648; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3650 = 7'h42 == io_i_rename_table_28 ? io_i_pregs_66 : _GEN_3649; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3651 = 7'h43 == io_i_rename_table_28 ? io_i_pregs_67 : _GEN_3650; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3652 = 7'h44 == io_i_rename_table_28 ? io_i_pregs_68 : _GEN_3651; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3653 = 7'h45 == io_i_rename_table_28 ? io_i_pregs_69 : _GEN_3652; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3654 = 7'h46 == io_i_rename_table_28 ? io_i_pregs_70 : _GEN_3653; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3655 = 7'h47 == io_i_rename_table_28 ? io_i_pregs_71 : _GEN_3654; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3656 = 7'h48 == io_i_rename_table_28 ? io_i_pregs_72 : _GEN_3655; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3657 = 7'h49 == io_i_rename_table_28 ? io_i_pregs_73 : _GEN_3656; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3658 = 7'h4a == io_i_rename_table_28 ? io_i_pregs_74 : _GEN_3657; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3659 = 7'h4b == io_i_rename_table_28 ? io_i_pregs_75 : _GEN_3658; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3660 = 7'h4c == io_i_rename_table_28 ? io_i_pregs_76 : _GEN_3659; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3661 = 7'h4d == io_i_rename_table_28 ? io_i_pregs_77 : _GEN_3660; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3662 = 7'h4e == io_i_rename_table_28 ? io_i_pregs_78 : _GEN_3661; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3663 = 7'h4f == io_i_rename_table_28 ? io_i_pregs_79 : _GEN_3662; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3664 = 7'h50 == io_i_rename_table_28 ? io_i_pregs_80 : _GEN_3663; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3665 = 7'h51 == io_i_rename_table_28 ? io_i_pregs_81 : _GEN_3664; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3666 = 7'h52 == io_i_rename_table_28 ? io_i_pregs_82 : _GEN_3665; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3667 = 7'h53 == io_i_rename_table_28 ? io_i_pregs_83 : _GEN_3666; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3668 = 7'h54 == io_i_rename_table_28 ? io_i_pregs_84 : _GEN_3667; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3669 = 7'h55 == io_i_rename_table_28 ? io_i_pregs_85 : _GEN_3668; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3670 = 7'h56 == io_i_rename_table_28 ? io_i_pregs_86 : _GEN_3669; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3671 = 7'h57 == io_i_rename_table_28 ? io_i_pregs_87 : _GEN_3670; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3672 = 7'h58 == io_i_rename_table_28 ? io_i_pregs_88 : _GEN_3671; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3673 = 7'h59 == io_i_rename_table_28 ? io_i_pregs_89 : _GEN_3672; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3674 = 7'h5a == io_i_rename_table_28 ? io_i_pregs_90 : _GEN_3673; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3675 = 7'h5b == io_i_rename_table_28 ? io_i_pregs_91 : _GEN_3674; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3676 = 7'h5c == io_i_rename_table_28 ? io_i_pregs_92 : _GEN_3675; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3677 = 7'h5d == io_i_rename_table_28 ? io_i_pregs_93 : _GEN_3676; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3678 = 7'h5e == io_i_rename_table_28 ? io_i_pregs_94 : _GEN_3677; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3679 = 7'h5f == io_i_rename_table_28 ? io_i_pregs_95 : _GEN_3678; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3680 = 7'h60 == io_i_rename_table_28 ? io_i_pregs_96 : _GEN_3679; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3681 = 7'h61 == io_i_rename_table_28 ? io_i_pregs_97 : _GEN_3680; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3682 = 7'h62 == io_i_rename_table_28 ? io_i_pregs_98 : _GEN_3681; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3683 = 7'h63 == io_i_rename_table_28 ? io_i_pregs_99 : _GEN_3682; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3684 = 7'h64 == io_i_rename_table_28 ? io_i_pregs_100 : _GEN_3683; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3685 = 7'h65 == io_i_rename_table_28 ? io_i_pregs_101 : _GEN_3684; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3686 = 7'h66 == io_i_rename_table_28 ? io_i_pregs_102 : _GEN_3685; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3687 = 7'h67 == io_i_rename_table_28 ? io_i_pregs_103 : _GEN_3686; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3688 = 7'h68 == io_i_rename_table_28 ? io_i_pregs_104 : _GEN_3687; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3689 = 7'h69 == io_i_rename_table_28 ? io_i_pregs_105 : _GEN_3688; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3690 = 7'h6a == io_i_rename_table_28 ? io_i_pregs_106 : _GEN_3689; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3691 = 7'h6b == io_i_rename_table_28 ? io_i_pregs_107 : _GEN_3690; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3692 = 7'h6c == io_i_rename_table_28 ? io_i_pregs_108 : _GEN_3691; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3693 = 7'h6d == io_i_rename_table_28 ? io_i_pregs_109 : _GEN_3692; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3694 = 7'h6e == io_i_rename_table_28 ? io_i_pregs_110 : _GEN_3693; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3695 = 7'h6f == io_i_rename_table_28 ? io_i_pregs_111 : _GEN_3694; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3696 = 7'h70 == io_i_rename_table_28 ? io_i_pregs_112 : _GEN_3695; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3697 = 7'h71 == io_i_rename_table_28 ? io_i_pregs_113 : _GEN_3696; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3698 = 7'h72 == io_i_rename_table_28 ? io_i_pregs_114 : _GEN_3697; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3699 = 7'h73 == io_i_rename_table_28 ? io_i_pregs_115 : _GEN_3698; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3700 = 7'h74 == io_i_rename_table_28 ? io_i_pregs_116 : _GEN_3699; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3701 = 7'h75 == io_i_rename_table_28 ? io_i_pregs_117 : _GEN_3700; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3702 = 7'h76 == io_i_rename_table_28 ? io_i_pregs_118 : _GEN_3701; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3703 = 7'h77 == io_i_rename_table_28 ? io_i_pregs_119 : _GEN_3702; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3704 = 7'h78 == io_i_rename_table_28 ? io_i_pregs_120 : _GEN_3703; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3705 = 7'h79 == io_i_rename_table_28 ? io_i_pregs_121 : _GEN_3704; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3706 = 7'h7a == io_i_rename_table_28 ? io_i_pregs_122 : _GEN_3705; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3707 = 7'h7b == io_i_rename_table_28 ? io_i_pregs_123 : _GEN_3706; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3708 = 7'h7c == io_i_rename_table_28 ? io_i_pregs_124 : _GEN_3707; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3709 = 7'h7d == io_i_rename_table_28 ? io_i_pregs_125 : _GEN_3708; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3710 = 7'h7e == io_i_rename_table_28 ? io_i_pregs_126 : _GEN_3709; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3713 = 7'h1 == io_i_rename_table_29 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3714 = 7'h2 == io_i_rename_table_29 ? io_i_pregs_2 : _GEN_3713; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3715 = 7'h3 == io_i_rename_table_29 ? io_i_pregs_3 : _GEN_3714; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3716 = 7'h4 == io_i_rename_table_29 ? io_i_pregs_4 : _GEN_3715; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3717 = 7'h5 == io_i_rename_table_29 ? io_i_pregs_5 : _GEN_3716; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3718 = 7'h6 == io_i_rename_table_29 ? io_i_pregs_6 : _GEN_3717; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3719 = 7'h7 == io_i_rename_table_29 ? io_i_pregs_7 : _GEN_3718; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3720 = 7'h8 == io_i_rename_table_29 ? io_i_pregs_8 : _GEN_3719; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3721 = 7'h9 == io_i_rename_table_29 ? io_i_pregs_9 : _GEN_3720; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3722 = 7'ha == io_i_rename_table_29 ? io_i_pregs_10 : _GEN_3721; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3723 = 7'hb == io_i_rename_table_29 ? io_i_pregs_11 : _GEN_3722; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3724 = 7'hc == io_i_rename_table_29 ? io_i_pregs_12 : _GEN_3723; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3725 = 7'hd == io_i_rename_table_29 ? io_i_pregs_13 : _GEN_3724; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3726 = 7'he == io_i_rename_table_29 ? io_i_pregs_14 : _GEN_3725; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3727 = 7'hf == io_i_rename_table_29 ? io_i_pregs_15 : _GEN_3726; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3728 = 7'h10 == io_i_rename_table_29 ? io_i_pregs_16 : _GEN_3727; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3729 = 7'h11 == io_i_rename_table_29 ? io_i_pregs_17 : _GEN_3728; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3730 = 7'h12 == io_i_rename_table_29 ? io_i_pregs_18 : _GEN_3729; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3731 = 7'h13 == io_i_rename_table_29 ? io_i_pregs_19 : _GEN_3730; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3732 = 7'h14 == io_i_rename_table_29 ? io_i_pregs_20 : _GEN_3731; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3733 = 7'h15 == io_i_rename_table_29 ? io_i_pregs_21 : _GEN_3732; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3734 = 7'h16 == io_i_rename_table_29 ? io_i_pregs_22 : _GEN_3733; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3735 = 7'h17 == io_i_rename_table_29 ? io_i_pregs_23 : _GEN_3734; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3736 = 7'h18 == io_i_rename_table_29 ? io_i_pregs_24 : _GEN_3735; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3737 = 7'h19 == io_i_rename_table_29 ? io_i_pregs_25 : _GEN_3736; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3738 = 7'h1a == io_i_rename_table_29 ? io_i_pregs_26 : _GEN_3737; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3739 = 7'h1b == io_i_rename_table_29 ? io_i_pregs_27 : _GEN_3738; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3740 = 7'h1c == io_i_rename_table_29 ? io_i_pregs_28 : _GEN_3739; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3741 = 7'h1d == io_i_rename_table_29 ? io_i_pregs_29 : _GEN_3740; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3742 = 7'h1e == io_i_rename_table_29 ? io_i_pregs_30 : _GEN_3741; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3743 = 7'h1f == io_i_rename_table_29 ? io_i_pregs_31 : _GEN_3742; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3744 = 7'h20 == io_i_rename_table_29 ? io_i_pregs_32 : _GEN_3743; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3745 = 7'h21 == io_i_rename_table_29 ? io_i_pregs_33 : _GEN_3744; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3746 = 7'h22 == io_i_rename_table_29 ? io_i_pregs_34 : _GEN_3745; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3747 = 7'h23 == io_i_rename_table_29 ? io_i_pregs_35 : _GEN_3746; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3748 = 7'h24 == io_i_rename_table_29 ? io_i_pregs_36 : _GEN_3747; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3749 = 7'h25 == io_i_rename_table_29 ? io_i_pregs_37 : _GEN_3748; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3750 = 7'h26 == io_i_rename_table_29 ? io_i_pregs_38 : _GEN_3749; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3751 = 7'h27 == io_i_rename_table_29 ? io_i_pregs_39 : _GEN_3750; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3752 = 7'h28 == io_i_rename_table_29 ? io_i_pregs_40 : _GEN_3751; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3753 = 7'h29 == io_i_rename_table_29 ? io_i_pregs_41 : _GEN_3752; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3754 = 7'h2a == io_i_rename_table_29 ? io_i_pregs_42 : _GEN_3753; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3755 = 7'h2b == io_i_rename_table_29 ? io_i_pregs_43 : _GEN_3754; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3756 = 7'h2c == io_i_rename_table_29 ? io_i_pregs_44 : _GEN_3755; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3757 = 7'h2d == io_i_rename_table_29 ? io_i_pregs_45 : _GEN_3756; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3758 = 7'h2e == io_i_rename_table_29 ? io_i_pregs_46 : _GEN_3757; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3759 = 7'h2f == io_i_rename_table_29 ? io_i_pregs_47 : _GEN_3758; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3760 = 7'h30 == io_i_rename_table_29 ? io_i_pregs_48 : _GEN_3759; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3761 = 7'h31 == io_i_rename_table_29 ? io_i_pregs_49 : _GEN_3760; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3762 = 7'h32 == io_i_rename_table_29 ? io_i_pregs_50 : _GEN_3761; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3763 = 7'h33 == io_i_rename_table_29 ? io_i_pregs_51 : _GEN_3762; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3764 = 7'h34 == io_i_rename_table_29 ? io_i_pregs_52 : _GEN_3763; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3765 = 7'h35 == io_i_rename_table_29 ? io_i_pregs_53 : _GEN_3764; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3766 = 7'h36 == io_i_rename_table_29 ? io_i_pregs_54 : _GEN_3765; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3767 = 7'h37 == io_i_rename_table_29 ? io_i_pregs_55 : _GEN_3766; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3768 = 7'h38 == io_i_rename_table_29 ? io_i_pregs_56 : _GEN_3767; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3769 = 7'h39 == io_i_rename_table_29 ? io_i_pregs_57 : _GEN_3768; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3770 = 7'h3a == io_i_rename_table_29 ? io_i_pregs_58 : _GEN_3769; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3771 = 7'h3b == io_i_rename_table_29 ? io_i_pregs_59 : _GEN_3770; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3772 = 7'h3c == io_i_rename_table_29 ? io_i_pregs_60 : _GEN_3771; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3773 = 7'h3d == io_i_rename_table_29 ? io_i_pregs_61 : _GEN_3772; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3774 = 7'h3e == io_i_rename_table_29 ? io_i_pregs_62 : _GEN_3773; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3775 = 7'h3f == io_i_rename_table_29 ? io_i_pregs_63 : _GEN_3774; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3776 = 7'h40 == io_i_rename_table_29 ? io_i_pregs_64 : _GEN_3775; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3777 = 7'h41 == io_i_rename_table_29 ? io_i_pregs_65 : _GEN_3776; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3778 = 7'h42 == io_i_rename_table_29 ? io_i_pregs_66 : _GEN_3777; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3779 = 7'h43 == io_i_rename_table_29 ? io_i_pregs_67 : _GEN_3778; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3780 = 7'h44 == io_i_rename_table_29 ? io_i_pregs_68 : _GEN_3779; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3781 = 7'h45 == io_i_rename_table_29 ? io_i_pregs_69 : _GEN_3780; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3782 = 7'h46 == io_i_rename_table_29 ? io_i_pregs_70 : _GEN_3781; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3783 = 7'h47 == io_i_rename_table_29 ? io_i_pregs_71 : _GEN_3782; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3784 = 7'h48 == io_i_rename_table_29 ? io_i_pregs_72 : _GEN_3783; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3785 = 7'h49 == io_i_rename_table_29 ? io_i_pregs_73 : _GEN_3784; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3786 = 7'h4a == io_i_rename_table_29 ? io_i_pregs_74 : _GEN_3785; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3787 = 7'h4b == io_i_rename_table_29 ? io_i_pregs_75 : _GEN_3786; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3788 = 7'h4c == io_i_rename_table_29 ? io_i_pregs_76 : _GEN_3787; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3789 = 7'h4d == io_i_rename_table_29 ? io_i_pregs_77 : _GEN_3788; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3790 = 7'h4e == io_i_rename_table_29 ? io_i_pregs_78 : _GEN_3789; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3791 = 7'h4f == io_i_rename_table_29 ? io_i_pregs_79 : _GEN_3790; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3792 = 7'h50 == io_i_rename_table_29 ? io_i_pregs_80 : _GEN_3791; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3793 = 7'h51 == io_i_rename_table_29 ? io_i_pregs_81 : _GEN_3792; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3794 = 7'h52 == io_i_rename_table_29 ? io_i_pregs_82 : _GEN_3793; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3795 = 7'h53 == io_i_rename_table_29 ? io_i_pregs_83 : _GEN_3794; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3796 = 7'h54 == io_i_rename_table_29 ? io_i_pregs_84 : _GEN_3795; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3797 = 7'h55 == io_i_rename_table_29 ? io_i_pregs_85 : _GEN_3796; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3798 = 7'h56 == io_i_rename_table_29 ? io_i_pregs_86 : _GEN_3797; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3799 = 7'h57 == io_i_rename_table_29 ? io_i_pregs_87 : _GEN_3798; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3800 = 7'h58 == io_i_rename_table_29 ? io_i_pregs_88 : _GEN_3799; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3801 = 7'h59 == io_i_rename_table_29 ? io_i_pregs_89 : _GEN_3800; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3802 = 7'h5a == io_i_rename_table_29 ? io_i_pregs_90 : _GEN_3801; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3803 = 7'h5b == io_i_rename_table_29 ? io_i_pregs_91 : _GEN_3802; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3804 = 7'h5c == io_i_rename_table_29 ? io_i_pregs_92 : _GEN_3803; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3805 = 7'h5d == io_i_rename_table_29 ? io_i_pregs_93 : _GEN_3804; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3806 = 7'h5e == io_i_rename_table_29 ? io_i_pregs_94 : _GEN_3805; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3807 = 7'h5f == io_i_rename_table_29 ? io_i_pregs_95 : _GEN_3806; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3808 = 7'h60 == io_i_rename_table_29 ? io_i_pregs_96 : _GEN_3807; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3809 = 7'h61 == io_i_rename_table_29 ? io_i_pregs_97 : _GEN_3808; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3810 = 7'h62 == io_i_rename_table_29 ? io_i_pregs_98 : _GEN_3809; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3811 = 7'h63 == io_i_rename_table_29 ? io_i_pregs_99 : _GEN_3810; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3812 = 7'h64 == io_i_rename_table_29 ? io_i_pregs_100 : _GEN_3811; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3813 = 7'h65 == io_i_rename_table_29 ? io_i_pregs_101 : _GEN_3812; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3814 = 7'h66 == io_i_rename_table_29 ? io_i_pregs_102 : _GEN_3813; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3815 = 7'h67 == io_i_rename_table_29 ? io_i_pregs_103 : _GEN_3814; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3816 = 7'h68 == io_i_rename_table_29 ? io_i_pregs_104 : _GEN_3815; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3817 = 7'h69 == io_i_rename_table_29 ? io_i_pregs_105 : _GEN_3816; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3818 = 7'h6a == io_i_rename_table_29 ? io_i_pregs_106 : _GEN_3817; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3819 = 7'h6b == io_i_rename_table_29 ? io_i_pregs_107 : _GEN_3818; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3820 = 7'h6c == io_i_rename_table_29 ? io_i_pregs_108 : _GEN_3819; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3821 = 7'h6d == io_i_rename_table_29 ? io_i_pregs_109 : _GEN_3820; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3822 = 7'h6e == io_i_rename_table_29 ? io_i_pregs_110 : _GEN_3821; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3823 = 7'h6f == io_i_rename_table_29 ? io_i_pregs_111 : _GEN_3822; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3824 = 7'h70 == io_i_rename_table_29 ? io_i_pregs_112 : _GEN_3823; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3825 = 7'h71 == io_i_rename_table_29 ? io_i_pregs_113 : _GEN_3824; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3826 = 7'h72 == io_i_rename_table_29 ? io_i_pregs_114 : _GEN_3825; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3827 = 7'h73 == io_i_rename_table_29 ? io_i_pregs_115 : _GEN_3826; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3828 = 7'h74 == io_i_rename_table_29 ? io_i_pregs_116 : _GEN_3827; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3829 = 7'h75 == io_i_rename_table_29 ? io_i_pregs_117 : _GEN_3828; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3830 = 7'h76 == io_i_rename_table_29 ? io_i_pregs_118 : _GEN_3829; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3831 = 7'h77 == io_i_rename_table_29 ? io_i_pregs_119 : _GEN_3830; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3832 = 7'h78 == io_i_rename_table_29 ? io_i_pregs_120 : _GEN_3831; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3833 = 7'h79 == io_i_rename_table_29 ? io_i_pregs_121 : _GEN_3832; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3834 = 7'h7a == io_i_rename_table_29 ? io_i_pregs_122 : _GEN_3833; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3835 = 7'h7b == io_i_rename_table_29 ? io_i_pregs_123 : _GEN_3834; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3836 = 7'h7c == io_i_rename_table_29 ? io_i_pregs_124 : _GEN_3835; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3837 = 7'h7d == io_i_rename_table_29 ? io_i_pregs_125 : _GEN_3836; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3838 = 7'h7e == io_i_rename_table_29 ? io_i_pregs_126 : _GEN_3837; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3841 = 7'h1 == io_i_rename_table_30 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3842 = 7'h2 == io_i_rename_table_30 ? io_i_pregs_2 : _GEN_3841; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3843 = 7'h3 == io_i_rename_table_30 ? io_i_pregs_3 : _GEN_3842; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3844 = 7'h4 == io_i_rename_table_30 ? io_i_pregs_4 : _GEN_3843; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3845 = 7'h5 == io_i_rename_table_30 ? io_i_pregs_5 : _GEN_3844; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3846 = 7'h6 == io_i_rename_table_30 ? io_i_pregs_6 : _GEN_3845; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3847 = 7'h7 == io_i_rename_table_30 ? io_i_pregs_7 : _GEN_3846; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3848 = 7'h8 == io_i_rename_table_30 ? io_i_pregs_8 : _GEN_3847; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3849 = 7'h9 == io_i_rename_table_30 ? io_i_pregs_9 : _GEN_3848; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3850 = 7'ha == io_i_rename_table_30 ? io_i_pregs_10 : _GEN_3849; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3851 = 7'hb == io_i_rename_table_30 ? io_i_pregs_11 : _GEN_3850; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3852 = 7'hc == io_i_rename_table_30 ? io_i_pregs_12 : _GEN_3851; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3853 = 7'hd == io_i_rename_table_30 ? io_i_pregs_13 : _GEN_3852; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3854 = 7'he == io_i_rename_table_30 ? io_i_pregs_14 : _GEN_3853; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3855 = 7'hf == io_i_rename_table_30 ? io_i_pregs_15 : _GEN_3854; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3856 = 7'h10 == io_i_rename_table_30 ? io_i_pregs_16 : _GEN_3855; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3857 = 7'h11 == io_i_rename_table_30 ? io_i_pregs_17 : _GEN_3856; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3858 = 7'h12 == io_i_rename_table_30 ? io_i_pregs_18 : _GEN_3857; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3859 = 7'h13 == io_i_rename_table_30 ? io_i_pregs_19 : _GEN_3858; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3860 = 7'h14 == io_i_rename_table_30 ? io_i_pregs_20 : _GEN_3859; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3861 = 7'h15 == io_i_rename_table_30 ? io_i_pregs_21 : _GEN_3860; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3862 = 7'h16 == io_i_rename_table_30 ? io_i_pregs_22 : _GEN_3861; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3863 = 7'h17 == io_i_rename_table_30 ? io_i_pregs_23 : _GEN_3862; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3864 = 7'h18 == io_i_rename_table_30 ? io_i_pregs_24 : _GEN_3863; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3865 = 7'h19 == io_i_rename_table_30 ? io_i_pregs_25 : _GEN_3864; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3866 = 7'h1a == io_i_rename_table_30 ? io_i_pregs_26 : _GEN_3865; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3867 = 7'h1b == io_i_rename_table_30 ? io_i_pregs_27 : _GEN_3866; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3868 = 7'h1c == io_i_rename_table_30 ? io_i_pregs_28 : _GEN_3867; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3869 = 7'h1d == io_i_rename_table_30 ? io_i_pregs_29 : _GEN_3868; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3870 = 7'h1e == io_i_rename_table_30 ? io_i_pregs_30 : _GEN_3869; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3871 = 7'h1f == io_i_rename_table_30 ? io_i_pregs_31 : _GEN_3870; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3872 = 7'h20 == io_i_rename_table_30 ? io_i_pregs_32 : _GEN_3871; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3873 = 7'h21 == io_i_rename_table_30 ? io_i_pregs_33 : _GEN_3872; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3874 = 7'h22 == io_i_rename_table_30 ? io_i_pregs_34 : _GEN_3873; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3875 = 7'h23 == io_i_rename_table_30 ? io_i_pregs_35 : _GEN_3874; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3876 = 7'h24 == io_i_rename_table_30 ? io_i_pregs_36 : _GEN_3875; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3877 = 7'h25 == io_i_rename_table_30 ? io_i_pregs_37 : _GEN_3876; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3878 = 7'h26 == io_i_rename_table_30 ? io_i_pregs_38 : _GEN_3877; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3879 = 7'h27 == io_i_rename_table_30 ? io_i_pregs_39 : _GEN_3878; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3880 = 7'h28 == io_i_rename_table_30 ? io_i_pregs_40 : _GEN_3879; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3881 = 7'h29 == io_i_rename_table_30 ? io_i_pregs_41 : _GEN_3880; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3882 = 7'h2a == io_i_rename_table_30 ? io_i_pregs_42 : _GEN_3881; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3883 = 7'h2b == io_i_rename_table_30 ? io_i_pregs_43 : _GEN_3882; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3884 = 7'h2c == io_i_rename_table_30 ? io_i_pregs_44 : _GEN_3883; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3885 = 7'h2d == io_i_rename_table_30 ? io_i_pregs_45 : _GEN_3884; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3886 = 7'h2e == io_i_rename_table_30 ? io_i_pregs_46 : _GEN_3885; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3887 = 7'h2f == io_i_rename_table_30 ? io_i_pregs_47 : _GEN_3886; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3888 = 7'h30 == io_i_rename_table_30 ? io_i_pregs_48 : _GEN_3887; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3889 = 7'h31 == io_i_rename_table_30 ? io_i_pregs_49 : _GEN_3888; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3890 = 7'h32 == io_i_rename_table_30 ? io_i_pregs_50 : _GEN_3889; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3891 = 7'h33 == io_i_rename_table_30 ? io_i_pregs_51 : _GEN_3890; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3892 = 7'h34 == io_i_rename_table_30 ? io_i_pregs_52 : _GEN_3891; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3893 = 7'h35 == io_i_rename_table_30 ? io_i_pregs_53 : _GEN_3892; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3894 = 7'h36 == io_i_rename_table_30 ? io_i_pregs_54 : _GEN_3893; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3895 = 7'h37 == io_i_rename_table_30 ? io_i_pregs_55 : _GEN_3894; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3896 = 7'h38 == io_i_rename_table_30 ? io_i_pregs_56 : _GEN_3895; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3897 = 7'h39 == io_i_rename_table_30 ? io_i_pregs_57 : _GEN_3896; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3898 = 7'h3a == io_i_rename_table_30 ? io_i_pregs_58 : _GEN_3897; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3899 = 7'h3b == io_i_rename_table_30 ? io_i_pregs_59 : _GEN_3898; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3900 = 7'h3c == io_i_rename_table_30 ? io_i_pregs_60 : _GEN_3899; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3901 = 7'h3d == io_i_rename_table_30 ? io_i_pregs_61 : _GEN_3900; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3902 = 7'h3e == io_i_rename_table_30 ? io_i_pregs_62 : _GEN_3901; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3903 = 7'h3f == io_i_rename_table_30 ? io_i_pregs_63 : _GEN_3902; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3904 = 7'h40 == io_i_rename_table_30 ? io_i_pregs_64 : _GEN_3903; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3905 = 7'h41 == io_i_rename_table_30 ? io_i_pregs_65 : _GEN_3904; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3906 = 7'h42 == io_i_rename_table_30 ? io_i_pregs_66 : _GEN_3905; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3907 = 7'h43 == io_i_rename_table_30 ? io_i_pregs_67 : _GEN_3906; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3908 = 7'h44 == io_i_rename_table_30 ? io_i_pregs_68 : _GEN_3907; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3909 = 7'h45 == io_i_rename_table_30 ? io_i_pregs_69 : _GEN_3908; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3910 = 7'h46 == io_i_rename_table_30 ? io_i_pregs_70 : _GEN_3909; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3911 = 7'h47 == io_i_rename_table_30 ? io_i_pregs_71 : _GEN_3910; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3912 = 7'h48 == io_i_rename_table_30 ? io_i_pregs_72 : _GEN_3911; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3913 = 7'h49 == io_i_rename_table_30 ? io_i_pregs_73 : _GEN_3912; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3914 = 7'h4a == io_i_rename_table_30 ? io_i_pregs_74 : _GEN_3913; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3915 = 7'h4b == io_i_rename_table_30 ? io_i_pregs_75 : _GEN_3914; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3916 = 7'h4c == io_i_rename_table_30 ? io_i_pregs_76 : _GEN_3915; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3917 = 7'h4d == io_i_rename_table_30 ? io_i_pregs_77 : _GEN_3916; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3918 = 7'h4e == io_i_rename_table_30 ? io_i_pregs_78 : _GEN_3917; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3919 = 7'h4f == io_i_rename_table_30 ? io_i_pregs_79 : _GEN_3918; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3920 = 7'h50 == io_i_rename_table_30 ? io_i_pregs_80 : _GEN_3919; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3921 = 7'h51 == io_i_rename_table_30 ? io_i_pregs_81 : _GEN_3920; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3922 = 7'h52 == io_i_rename_table_30 ? io_i_pregs_82 : _GEN_3921; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3923 = 7'h53 == io_i_rename_table_30 ? io_i_pregs_83 : _GEN_3922; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3924 = 7'h54 == io_i_rename_table_30 ? io_i_pregs_84 : _GEN_3923; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3925 = 7'h55 == io_i_rename_table_30 ? io_i_pregs_85 : _GEN_3924; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3926 = 7'h56 == io_i_rename_table_30 ? io_i_pregs_86 : _GEN_3925; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3927 = 7'h57 == io_i_rename_table_30 ? io_i_pregs_87 : _GEN_3926; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3928 = 7'h58 == io_i_rename_table_30 ? io_i_pregs_88 : _GEN_3927; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3929 = 7'h59 == io_i_rename_table_30 ? io_i_pregs_89 : _GEN_3928; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3930 = 7'h5a == io_i_rename_table_30 ? io_i_pregs_90 : _GEN_3929; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3931 = 7'h5b == io_i_rename_table_30 ? io_i_pregs_91 : _GEN_3930; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3932 = 7'h5c == io_i_rename_table_30 ? io_i_pregs_92 : _GEN_3931; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3933 = 7'h5d == io_i_rename_table_30 ? io_i_pregs_93 : _GEN_3932; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3934 = 7'h5e == io_i_rename_table_30 ? io_i_pregs_94 : _GEN_3933; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3935 = 7'h5f == io_i_rename_table_30 ? io_i_pregs_95 : _GEN_3934; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3936 = 7'h60 == io_i_rename_table_30 ? io_i_pregs_96 : _GEN_3935; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3937 = 7'h61 == io_i_rename_table_30 ? io_i_pregs_97 : _GEN_3936; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3938 = 7'h62 == io_i_rename_table_30 ? io_i_pregs_98 : _GEN_3937; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3939 = 7'h63 == io_i_rename_table_30 ? io_i_pregs_99 : _GEN_3938; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3940 = 7'h64 == io_i_rename_table_30 ? io_i_pregs_100 : _GEN_3939; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3941 = 7'h65 == io_i_rename_table_30 ? io_i_pregs_101 : _GEN_3940; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3942 = 7'h66 == io_i_rename_table_30 ? io_i_pregs_102 : _GEN_3941; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3943 = 7'h67 == io_i_rename_table_30 ? io_i_pregs_103 : _GEN_3942; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3944 = 7'h68 == io_i_rename_table_30 ? io_i_pregs_104 : _GEN_3943; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3945 = 7'h69 == io_i_rename_table_30 ? io_i_pregs_105 : _GEN_3944; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3946 = 7'h6a == io_i_rename_table_30 ? io_i_pregs_106 : _GEN_3945; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3947 = 7'h6b == io_i_rename_table_30 ? io_i_pregs_107 : _GEN_3946; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3948 = 7'h6c == io_i_rename_table_30 ? io_i_pregs_108 : _GEN_3947; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3949 = 7'h6d == io_i_rename_table_30 ? io_i_pregs_109 : _GEN_3948; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3950 = 7'h6e == io_i_rename_table_30 ? io_i_pregs_110 : _GEN_3949; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3951 = 7'h6f == io_i_rename_table_30 ? io_i_pregs_111 : _GEN_3950; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3952 = 7'h70 == io_i_rename_table_30 ? io_i_pregs_112 : _GEN_3951; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3953 = 7'h71 == io_i_rename_table_30 ? io_i_pregs_113 : _GEN_3952; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3954 = 7'h72 == io_i_rename_table_30 ? io_i_pregs_114 : _GEN_3953; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3955 = 7'h73 == io_i_rename_table_30 ? io_i_pregs_115 : _GEN_3954; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3956 = 7'h74 == io_i_rename_table_30 ? io_i_pregs_116 : _GEN_3955; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3957 = 7'h75 == io_i_rename_table_30 ? io_i_pregs_117 : _GEN_3956; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3958 = 7'h76 == io_i_rename_table_30 ? io_i_pregs_118 : _GEN_3957; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3959 = 7'h77 == io_i_rename_table_30 ? io_i_pregs_119 : _GEN_3958; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3960 = 7'h78 == io_i_rename_table_30 ? io_i_pregs_120 : _GEN_3959; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3961 = 7'h79 == io_i_rename_table_30 ? io_i_pregs_121 : _GEN_3960; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3962 = 7'h7a == io_i_rename_table_30 ? io_i_pregs_122 : _GEN_3961; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3963 = 7'h7b == io_i_rename_table_30 ? io_i_pregs_123 : _GEN_3962; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3964 = 7'h7c == io_i_rename_table_30 ? io_i_pregs_124 : _GEN_3963; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3965 = 7'h7d == io_i_rename_table_30 ? io_i_pregs_125 : _GEN_3964; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3966 = 7'h7e == io_i_rename_table_30 ? io_i_pregs_126 : _GEN_3965; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3969 = 7'h1 == io_i_rename_table_31 ? io_i_pregs_1 : io_i_pregs_0; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3970 = 7'h2 == io_i_rename_table_31 ? io_i_pregs_2 : _GEN_3969; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3971 = 7'h3 == io_i_rename_table_31 ? io_i_pregs_3 : _GEN_3970; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3972 = 7'h4 == io_i_rename_table_31 ? io_i_pregs_4 : _GEN_3971; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3973 = 7'h5 == io_i_rename_table_31 ? io_i_pregs_5 : _GEN_3972; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3974 = 7'h6 == io_i_rename_table_31 ? io_i_pregs_6 : _GEN_3973; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3975 = 7'h7 == io_i_rename_table_31 ? io_i_pregs_7 : _GEN_3974; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3976 = 7'h8 == io_i_rename_table_31 ? io_i_pregs_8 : _GEN_3975; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3977 = 7'h9 == io_i_rename_table_31 ? io_i_pregs_9 : _GEN_3976; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3978 = 7'ha == io_i_rename_table_31 ? io_i_pregs_10 : _GEN_3977; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3979 = 7'hb == io_i_rename_table_31 ? io_i_pregs_11 : _GEN_3978; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3980 = 7'hc == io_i_rename_table_31 ? io_i_pregs_12 : _GEN_3979; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3981 = 7'hd == io_i_rename_table_31 ? io_i_pregs_13 : _GEN_3980; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3982 = 7'he == io_i_rename_table_31 ? io_i_pregs_14 : _GEN_3981; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3983 = 7'hf == io_i_rename_table_31 ? io_i_pregs_15 : _GEN_3982; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3984 = 7'h10 == io_i_rename_table_31 ? io_i_pregs_16 : _GEN_3983; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3985 = 7'h11 == io_i_rename_table_31 ? io_i_pregs_17 : _GEN_3984; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3986 = 7'h12 == io_i_rename_table_31 ? io_i_pregs_18 : _GEN_3985; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3987 = 7'h13 == io_i_rename_table_31 ? io_i_pregs_19 : _GEN_3986; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3988 = 7'h14 == io_i_rename_table_31 ? io_i_pregs_20 : _GEN_3987; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3989 = 7'h15 == io_i_rename_table_31 ? io_i_pregs_21 : _GEN_3988; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3990 = 7'h16 == io_i_rename_table_31 ? io_i_pregs_22 : _GEN_3989; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3991 = 7'h17 == io_i_rename_table_31 ? io_i_pregs_23 : _GEN_3990; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3992 = 7'h18 == io_i_rename_table_31 ? io_i_pregs_24 : _GEN_3991; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3993 = 7'h19 == io_i_rename_table_31 ? io_i_pregs_25 : _GEN_3992; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3994 = 7'h1a == io_i_rename_table_31 ? io_i_pregs_26 : _GEN_3993; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3995 = 7'h1b == io_i_rename_table_31 ? io_i_pregs_27 : _GEN_3994; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3996 = 7'h1c == io_i_rename_table_31 ? io_i_pregs_28 : _GEN_3995; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3997 = 7'h1d == io_i_rename_table_31 ? io_i_pregs_29 : _GEN_3996; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3998 = 7'h1e == io_i_rename_table_31 ? io_i_pregs_30 : _GEN_3997; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_3999 = 7'h1f == io_i_rename_table_31 ? io_i_pregs_31 : _GEN_3998; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4000 = 7'h20 == io_i_rename_table_31 ? io_i_pregs_32 : _GEN_3999; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4001 = 7'h21 == io_i_rename_table_31 ? io_i_pregs_33 : _GEN_4000; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4002 = 7'h22 == io_i_rename_table_31 ? io_i_pregs_34 : _GEN_4001; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4003 = 7'h23 == io_i_rename_table_31 ? io_i_pregs_35 : _GEN_4002; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4004 = 7'h24 == io_i_rename_table_31 ? io_i_pregs_36 : _GEN_4003; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4005 = 7'h25 == io_i_rename_table_31 ? io_i_pregs_37 : _GEN_4004; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4006 = 7'h26 == io_i_rename_table_31 ? io_i_pregs_38 : _GEN_4005; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4007 = 7'h27 == io_i_rename_table_31 ? io_i_pregs_39 : _GEN_4006; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4008 = 7'h28 == io_i_rename_table_31 ? io_i_pregs_40 : _GEN_4007; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4009 = 7'h29 == io_i_rename_table_31 ? io_i_pregs_41 : _GEN_4008; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4010 = 7'h2a == io_i_rename_table_31 ? io_i_pregs_42 : _GEN_4009; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4011 = 7'h2b == io_i_rename_table_31 ? io_i_pregs_43 : _GEN_4010; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4012 = 7'h2c == io_i_rename_table_31 ? io_i_pregs_44 : _GEN_4011; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4013 = 7'h2d == io_i_rename_table_31 ? io_i_pregs_45 : _GEN_4012; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4014 = 7'h2e == io_i_rename_table_31 ? io_i_pregs_46 : _GEN_4013; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4015 = 7'h2f == io_i_rename_table_31 ? io_i_pregs_47 : _GEN_4014; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4016 = 7'h30 == io_i_rename_table_31 ? io_i_pregs_48 : _GEN_4015; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4017 = 7'h31 == io_i_rename_table_31 ? io_i_pregs_49 : _GEN_4016; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4018 = 7'h32 == io_i_rename_table_31 ? io_i_pregs_50 : _GEN_4017; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4019 = 7'h33 == io_i_rename_table_31 ? io_i_pregs_51 : _GEN_4018; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4020 = 7'h34 == io_i_rename_table_31 ? io_i_pregs_52 : _GEN_4019; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4021 = 7'h35 == io_i_rename_table_31 ? io_i_pregs_53 : _GEN_4020; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4022 = 7'h36 == io_i_rename_table_31 ? io_i_pregs_54 : _GEN_4021; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4023 = 7'h37 == io_i_rename_table_31 ? io_i_pregs_55 : _GEN_4022; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4024 = 7'h38 == io_i_rename_table_31 ? io_i_pregs_56 : _GEN_4023; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4025 = 7'h39 == io_i_rename_table_31 ? io_i_pregs_57 : _GEN_4024; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4026 = 7'h3a == io_i_rename_table_31 ? io_i_pregs_58 : _GEN_4025; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4027 = 7'h3b == io_i_rename_table_31 ? io_i_pregs_59 : _GEN_4026; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4028 = 7'h3c == io_i_rename_table_31 ? io_i_pregs_60 : _GEN_4027; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4029 = 7'h3d == io_i_rename_table_31 ? io_i_pregs_61 : _GEN_4028; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4030 = 7'h3e == io_i_rename_table_31 ? io_i_pregs_62 : _GEN_4029; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4031 = 7'h3f == io_i_rename_table_31 ? io_i_pregs_63 : _GEN_4030; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4032 = 7'h40 == io_i_rename_table_31 ? io_i_pregs_64 : _GEN_4031; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4033 = 7'h41 == io_i_rename_table_31 ? io_i_pregs_65 : _GEN_4032; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4034 = 7'h42 == io_i_rename_table_31 ? io_i_pregs_66 : _GEN_4033; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4035 = 7'h43 == io_i_rename_table_31 ? io_i_pregs_67 : _GEN_4034; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4036 = 7'h44 == io_i_rename_table_31 ? io_i_pregs_68 : _GEN_4035; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4037 = 7'h45 == io_i_rename_table_31 ? io_i_pregs_69 : _GEN_4036; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4038 = 7'h46 == io_i_rename_table_31 ? io_i_pregs_70 : _GEN_4037; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4039 = 7'h47 == io_i_rename_table_31 ? io_i_pregs_71 : _GEN_4038; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4040 = 7'h48 == io_i_rename_table_31 ? io_i_pregs_72 : _GEN_4039; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4041 = 7'h49 == io_i_rename_table_31 ? io_i_pregs_73 : _GEN_4040; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4042 = 7'h4a == io_i_rename_table_31 ? io_i_pregs_74 : _GEN_4041; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4043 = 7'h4b == io_i_rename_table_31 ? io_i_pregs_75 : _GEN_4042; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4044 = 7'h4c == io_i_rename_table_31 ? io_i_pregs_76 : _GEN_4043; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4045 = 7'h4d == io_i_rename_table_31 ? io_i_pregs_77 : _GEN_4044; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4046 = 7'h4e == io_i_rename_table_31 ? io_i_pregs_78 : _GEN_4045; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4047 = 7'h4f == io_i_rename_table_31 ? io_i_pregs_79 : _GEN_4046; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4048 = 7'h50 == io_i_rename_table_31 ? io_i_pregs_80 : _GEN_4047; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4049 = 7'h51 == io_i_rename_table_31 ? io_i_pregs_81 : _GEN_4048; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4050 = 7'h52 == io_i_rename_table_31 ? io_i_pregs_82 : _GEN_4049; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4051 = 7'h53 == io_i_rename_table_31 ? io_i_pregs_83 : _GEN_4050; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4052 = 7'h54 == io_i_rename_table_31 ? io_i_pregs_84 : _GEN_4051; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4053 = 7'h55 == io_i_rename_table_31 ? io_i_pregs_85 : _GEN_4052; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4054 = 7'h56 == io_i_rename_table_31 ? io_i_pregs_86 : _GEN_4053; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4055 = 7'h57 == io_i_rename_table_31 ? io_i_pregs_87 : _GEN_4054; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4056 = 7'h58 == io_i_rename_table_31 ? io_i_pregs_88 : _GEN_4055; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4057 = 7'h59 == io_i_rename_table_31 ? io_i_pregs_89 : _GEN_4056; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4058 = 7'h5a == io_i_rename_table_31 ? io_i_pregs_90 : _GEN_4057; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4059 = 7'h5b == io_i_rename_table_31 ? io_i_pregs_91 : _GEN_4058; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4060 = 7'h5c == io_i_rename_table_31 ? io_i_pregs_92 : _GEN_4059; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4061 = 7'h5d == io_i_rename_table_31 ? io_i_pregs_93 : _GEN_4060; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4062 = 7'h5e == io_i_rename_table_31 ? io_i_pregs_94 : _GEN_4061; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4063 = 7'h5f == io_i_rename_table_31 ? io_i_pregs_95 : _GEN_4062; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4064 = 7'h60 == io_i_rename_table_31 ? io_i_pregs_96 : _GEN_4063; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4065 = 7'h61 == io_i_rename_table_31 ? io_i_pregs_97 : _GEN_4064; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4066 = 7'h62 == io_i_rename_table_31 ? io_i_pregs_98 : _GEN_4065; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4067 = 7'h63 == io_i_rename_table_31 ? io_i_pregs_99 : _GEN_4066; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4068 = 7'h64 == io_i_rename_table_31 ? io_i_pregs_100 : _GEN_4067; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4069 = 7'h65 == io_i_rename_table_31 ? io_i_pregs_101 : _GEN_4068; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4070 = 7'h66 == io_i_rename_table_31 ? io_i_pregs_102 : _GEN_4069; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4071 = 7'h67 == io_i_rename_table_31 ? io_i_pregs_103 : _GEN_4070; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4072 = 7'h68 == io_i_rename_table_31 ? io_i_pregs_104 : _GEN_4071; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4073 = 7'h69 == io_i_rename_table_31 ? io_i_pregs_105 : _GEN_4072; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4074 = 7'h6a == io_i_rename_table_31 ? io_i_pregs_106 : _GEN_4073; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4075 = 7'h6b == io_i_rename_table_31 ? io_i_pregs_107 : _GEN_4074; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4076 = 7'h6c == io_i_rename_table_31 ? io_i_pregs_108 : _GEN_4075; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4077 = 7'h6d == io_i_rename_table_31 ? io_i_pregs_109 : _GEN_4076; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4078 = 7'h6e == io_i_rename_table_31 ? io_i_pregs_110 : _GEN_4077; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4079 = 7'h6f == io_i_rename_table_31 ? io_i_pregs_111 : _GEN_4078; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4080 = 7'h70 == io_i_rename_table_31 ? io_i_pregs_112 : _GEN_4079; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4081 = 7'h71 == io_i_rename_table_31 ? io_i_pregs_113 : _GEN_4080; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4082 = 7'h72 == io_i_rename_table_31 ? io_i_pregs_114 : _GEN_4081; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4083 = 7'h73 == io_i_rename_table_31 ? io_i_pregs_115 : _GEN_4082; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4084 = 7'h74 == io_i_rename_table_31 ? io_i_pregs_116 : _GEN_4083; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4085 = 7'h75 == io_i_rename_table_31 ? io_i_pregs_117 : _GEN_4084; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4086 = 7'h76 == io_i_rename_table_31 ? io_i_pregs_118 : _GEN_4085; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4087 = 7'h77 == io_i_rename_table_31 ? io_i_pregs_119 : _GEN_4086; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4088 = 7'h78 == io_i_rename_table_31 ? io_i_pregs_120 : _GEN_4087; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4089 = 7'h79 == io_i_rename_table_31 ? io_i_pregs_121 : _GEN_4088; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4090 = 7'h7a == io_i_rename_table_31 ? io_i_pregs_122 : _GEN_4089; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4091 = 7'h7b == io_i_rename_table_31 ? io_i_pregs_123 : _GEN_4090; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4092 = 7'h7c == io_i_rename_table_31 ? io_i_pregs_124 : _GEN_4091; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4093 = 7'h7d == io_i_rename_table_31 ? io_i_pregs_125 : _GEN_4092; // @[arch_regfile.scala 21:{27,27}]
  wire [63:0] _GEN_4094 = 7'h7e == io_i_rename_table_31 ? io_i_pregs_126 : _GEN_4093; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_0 = 7'h7f == io_i_rename_table_0 ? io_i_pregs_127 : _GEN_126; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_1 = 7'h7f == io_i_rename_table_1 ? io_i_pregs_127 : _GEN_254; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_2 = 7'h7f == io_i_rename_table_2 ? io_i_pregs_127 : _GEN_382; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_3 = 7'h7f == io_i_rename_table_3 ? io_i_pregs_127 : _GEN_510; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_4 = 7'h7f == io_i_rename_table_4 ? io_i_pregs_127 : _GEN_638; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_5 = 7'h7f == io_i_rename_table_5 ? io_i_pregs_127 : _GEN_766; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_6 = 7'h7f == io_i_rename_table_6 ? io_i_pregs_127 : _GEN_894; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_7 = 7'h7f == io_i_rename_table_7 ? io_i_pregs_127 : _GEN_1022; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_8 = 7'h7f == io_i_rename_table_8 ? io_i_pregs_127 : _GEN_1150; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_9 = 7'h7f == io_i_rename_table_9 ? io_i_pregs_127 : _GEN_1278; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_10 = 7'h7f == io_i_rename_table_10 ? io_i_pregs_127 : _GEN_1406; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_11 = 7'h7f == io_i_rename_table_11 ? io_i_pregs_127 : _GEN_1534; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_12 = 7'h7f == io_i_rename_table_12 ? io_i_pregs_127 : _GEN_1662; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_13 = 7'h7f == io_i_rename_table_13 ? io_i_pregs_127 : _GEN_1790; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_14 = 7'h7f == io_i_rename_table_14 ? io_i_pregs_127 : _GEN_1918; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_15 = 7'h7f == io_i_rename_table_15 ? io_i_pregs_127 : _GEN_2046; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_16 = 7'h7f == io_i_rename_table_16 ? io_i_pregs_127 : _GEN_2174; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_17 = 7'h7f == io_i_rename_table_17 ? io_i_pregs_127 : _GEN_2302; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_18 = 7'h7f == io_i_rename_table_18 ? io_i_pregs_127 : _GEN_2430; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_19 = 7'h7f == io_i_rename_table_19 ? io_i_pregs_127 : _GEN_2558; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_20 = 7'h7f == io_i_rename_table_20 ? io_i_pregs_127 : _GEN_2686; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_21 = 7'h7f == io_i_rename_table_21 ? io_i_pregs_127 : _GEN_2814; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_22 = 7'h7f == io_i_rename_table_22 ? io_i_pregs_127 : _GEN_2942; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_23 = 7'h7f == io_i_rename_table_23 ? io_i_pregs_127 : _GEN_3070; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_24 = 7'h7f == io_i_rename_table_24 ? io_i_pregs_127 : _GEN_3198; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_25 = 7'h7f == io_i_rename_table_25 ? io_i_pregs_127 : _GEN_3326; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_26 = 7'h7f == io_i_rename_table_26 ? io_i_pregs_127 : _GEN_3454; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_27 = 7'h7f == io_i_rename_table_27 ? io_i_pregs_127 : _GEN_3582; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_28 = 7'h7f == io_i_rename_table_28 ? io_i_pregs_127 : _GEN_3710; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_29 = 7'h7f == io_i_rename_table_29 ? io_i_pregs_127 : _GEN_3838; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_30 = 7'h7f == io_i_rename_table_30 ? io_i_pregs_127 : _GEN_3966; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_arch_regs_31 = 7'h7f == io_i_rename_table_31 ? io_i_pregs_127 : _GEN_4094; // @[arch_regfile.scala 21:{27,27}]
  assign io_o_csr_regs_0 = io_i_csrs_0; // @[arch_regfile.scala 24:26]
  assign io_o_csr_regs_1 = io_i_csrs_1; // @[arch_regfile.scala 24:26]
  assign io_o_csr_regs_2 = io_i_csrs_2; // @[arch_regfile.scala 24:26]
  assign io_o_csr_regs_3 = io_i_csrs_3; // @[arch_regfile.scala 24:26]
endmodule
